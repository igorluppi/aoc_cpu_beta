module hard_disk(write_clock, read_clock, reset, trilha, setor, data, dataOut, hdWrite, hdRead);

	parameter DATA_WIDTH = 32; // X bits
	
	parameter HD_SETORES_BITS = 10;
	
	localparam HD_TRILHAS_SIZE = 32;
	localparam HD_SETORES_SIZE = 2**HD_SETORES_BITS;
	localparam HD_SIZE = HD_TRILHAS_SIZE*HD_SETORES_SIZE;
	
	input [DATA_WIDTH-1:0] data;
	input [DATA_WIDTH-1:0] trilha;
	input [DATA_WIDTH-1:0] setor;
	input reset, hdWrite, hdRead, write_clock, read_clock;
	
	output [DATA_WIDTH-1:0] dataOut;
	
	reg [DATA_WIDTH-1:0] dataRead;
	reg [DATA_WIDTH-1:0] HD [HD_SIZE-1:0]; // HD_SIZE words of 32-bit memory
	
	
	initial 
	begin : INIT

	/*Tabela de Programas Distribuida*/
	/*Header File*/
	/**
	* HD[i_0] = ativo;
	* HD[i_1] = identificador;
	* HD[i_2] = tamanho;
	*/
	/*Header File 01*/
	HD[3072] = 32'd1;
	HD[3073] = 32'd1;
	HD[3074] = 32'd140;
	/*Header File 02*/
	HD[4096] = 32'd1;
	HD[4097] = 32'd2;
	HD[4098] = 32'd250;
	/*Header File 03*/
	HD[5120] = 32'd1;
	HD[5121] = 32'd3;
	HD[5122] = 32'd63;
	/*Header File 04*/
	HD[6144] = 32'd1;
	HD[6145] = 32'd4;
	HD[6146] = 32'd106;
	/*Header File 05*/
	HD[7168] = 32'd1;
	HD[7169] = 32'd5;
	HD[7170] = 32'd99;
	/*Header File 06*/
	HD[8192] = 32'd1;
	HD[8193] = 32'd6;
	HD[8194] = 32'd48;
	/*Header File 07*/
	HD[9216] = 32'd1;
	HD[9217] = 32'd7;
	HD[9218] = 32'd55;
	/*Header File 08*/
	HD[10240] = 32'd1;
	HD[10241] = 32'd8;
	HD[10242] = 32'd33;
	/*Header File 09*/
	HD[11264] = 32'd1;
	HD[11265] = 32'd9;
	HD[11266] = 32'd102;
	/*Header File 10*/
	HD[12288] = 32'd1;
	HD[12289] = 32'd10;
	HD[12290] = 32'd66;
	/*Header File 11*/
	HD[13312] = 32'd1;
	HD[13313] = 32'd11;
	HD[13314] = 32'd8;
	/*Header File 12*/
	HD[14336] = 32'd1;
	HD[14337] = 32'd12;
	HD[14338] = 32'd8;
	/*Header File 13*/
	HD[15360] = 32'd1;
	HD[15361] = 32'd13;
	HD[15362] = 32'd160;
	
	
	
	/*Sistema Operacional - Size:2925*/
	/* Parameters: <mem_offset = 0> <priority_system = true> <index_begin = -1> */
	HD[0] = 32'b000101_00000_00000_0000000000000000; // li $global 0
	HD[1] = 32'b000011_00000_10101_0000000000100001; // addi $fp $global 33
	HD[2] = 32'b001011_00000000000000101101101010; // jump main
	HD[3] = 32'b001111_10110_10111_0000000000000000; // push $ra / syscall_io
	HD[4] = 32'b00000000000000000000000000000000; // noop / _label4_
	HD[5] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[6] = 32'b000000_00010_11001_00000_00000_010000; // move 25 2
	HD[7] = 32'b000000_11010_00000_00000_00000_010100; // jr 26
	HD[8] = 32'b00000000000000000000000000000000; // noop / _label5_
	HD[9] = 32'b000000_11001_00010_00000_00000_010000; // move 2 25
	HD[10] = 32'b001010_00010_00000_0000000000000000; // out 2
	HD[11] = 32'b000000_11010_00000_00000_00000_010100; // jr 26
	HD[12] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[13] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[14] = 32'b001111_10110_10111_0000000000000000; // push $ra / retoma_execucao_so
	HD[15] = 32'b00000000000000000000000000000000; // noop / _label0_
	HD[16] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[17] = 32'b000010_00000_00010_0000000000010011; // sw 2 $global 19
	HD[18] = 32'b00000000000000000000000000000000; // noop / _label3_
	HD[19] = 32'b101011_00000000000000000000000000; // intr_off
	HD[20] = 32'b000001_00000_00010_0000000000000110; // lw 2 $global 6
	HD[21] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[22] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[23] = 32'b000111_00010_00000_0000000000000011; // beq 2 $zero _ElseBegin0_
	HD[24] = 32'b001011_00000000000000001111100111; // jump _label1_
	HD[25] = 32'b001011_00000000000000000000011111; // jump _IfExit0_
	HD[26] = 32'b000001_00000_00010_0000000000000110; // lw 2 $global 6 / _ElseBegin0_
	HD[27] = 32'b000101_00000_00011_0000000000000010; // li 3 2
	HD[28] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[29] = 32'b000111_00010_00000_0000000000000010; // beq 2 $zero _IfExit1_
	HD[30] = 32'b001011_00000000000000010010110010; // jump _label2_
	HD[31] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _IfExit1_ _IfExit0_
	HD[32] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[33] = 32'b001111_10110_10111_0000000000000000; // push $ra / sleep
	HD[34] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[35] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[36] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[37] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[38] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[39] = 32'b000111_00010_00000_0000000000000110; // beq 2 $zero _ElseBegin2_
	HD[40] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[41] = 32'b000101_00000_00011_0001100001101010; // li 3 6250
	HD[42] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[43] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[44] = 32'b001011_00000000000000000000110011; // jump _IfExit2_
	HD[45] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin2_
	HD[46] = 32'b000101_00000_00011_0000000000011001; // li 3 25
	HD[47] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[48] = 32'b000101_00000_00011_0000000000000100; // li 3 4
	HD[49] = 32'b000000_00010_00011_00010_00000_001000; // div 2 2 3
	HD[50] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[51] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2 / _IfExit2_ _WhileBegin0_
	HD[52] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[53] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[54] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _WhileExit0_
	HD[55] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[56] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[57] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[58] = 32'b001011_00000000000000000000110011; // jump _WhileBegin0_
	HD[59] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _WhileExit0_
	HD[60] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[61] = 32'b001111_10110_10111_0000000000000000; // push $ra / vetor_existe_valor
	HD[62] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[63] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[64] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3 / _WhileBegin1_
	HD[65] = 32'b000001_10101_00011_0000000000000001; // lw 3 $fp 1
	HD[66] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[67] = 32'b000111_00010_00000_0000000000010000; // beq 2 $zero _WhileExit1_
	HD[68] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[69] = 32'b000001_10101_00011_0000000000000011; // lw 3 $fp 3
	HD[70] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[71] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
	HD[72] = 32'b000001_10101_00011_0000000000000010; // lw 3 $fp 2
	HD[73] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[74] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _IfExit3_
	HD[75] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3
	HD[76] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[77] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[78] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[79] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3 / _IfExit3_
	HD[80] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[81] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[82] = 32'b001011_00000000000000000001000000; // jump _WhileBegin1_
	HD[83] = 32'b000101_00000_00010_0000000000000000; // li 2 0 / _WhileExit1_
	HD[84] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[85] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[86] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[87] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[88] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[89] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[90] = 32'b001111_10110_10111_0000000000000000; // push $ra / mod
	HD[91] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[92] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[93] = 32'b000001_10101_00100_0000000000000001; // lw 4 $fp 1
	HD[94] = 32'b000000_00011_00100_00011_00000_001000; // div 3 3 4
	HD[95] = 32'b000001_10101_00100_0000000000000001; // lw 4 $fp 1
	HD[96] = 32'b000000_00011_00100_00011_00000_000111; // mult 3 3 4
	HD[97] = 32'b000000_00010_00011_00010_00000_000110; // sub 2 2 3
	HD[98] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[99] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[100] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[101] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[102] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[103] = 32'b001111_10110_10111_0000000000000000; // push $ra / print_value
	HD[104] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[105] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[106] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[107] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[108] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[109] = 32'b101000_00000000000000000001011010; // jal mod
	HD[110] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[111] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[112] = 32'b000011_00010_00010_0000000000110000; // addi 2 2 48
	HD[113] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[114] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[115] = 32'b000101_00000_00011_0000000000010000; // li 3 16
	HD[116] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[117] = 32'b000001_10101_00011_0000000000000010; // lw 3 $fp 2
	HD[118] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[119] = 32'b000001_10101_00011_0000000000000011; // lw 3 $fp 3
	HD[120] = 32'b100111_00010_00011_00011_00000000000; // lcdwrite 2 3 3
	HD[121] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[122] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[123] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[124] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[125] = 32'b000111_00010_00000_0000000000001110; // beq 2 $zero _ElseBegin4_
	HD[126] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[127] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[128] = 32'b000000_00010_00011_00010_00000_001000; // div 2 2 3
	HD[129] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[130] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[131] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[132] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[133] = 32'b101000_00000000000000000001011010; // jal mod
	HD[134] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[135] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[136] = 32'b000011_00010_00010_0000000000110000; // addi 2 2 48
	HD[137] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[138] = 32'b001011_00000000000000000010001101; // jump _IfExit4_
	HD[139] = 32'b000101_00000_00010_0000000000100000; // li 2 32 / _ElseBegin4_
	HD[140] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[141] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _IfExit4_
	HD[142] = 32'b000101_00000_00011_0000000000010000; // li 3 16
	HD[143] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[144] = 32'b000001_10101_00011_0000000000000010; // lw 3 $fp 2
	HD[145] = 32'b000100_00011_00011_0000000000000001; // subi 3 3 1
	HD[146] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[147] = 32'b000001_10101_00011_0000000000000011; // lw 3 $fp 3
	HD[148] = 32'b100111_00010_00011_00011_00000000000; // lcdwrite 2 3 3
	HD[149] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[150] = 32'b000101_00000_00011_0000000001100100; // li 3 100
	HD[151] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[152] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[153] = 32'b000111_00010_00000_0000000000001110; // beq 2 $zero _ElseBegin5_
	HD[154] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[155] = 32'b000101_00000_00011_0000000001100100; // li 3 100
	HD[156] = 32'b000000_00010_00011_00010_00000_001000; // div 2 2 3
	HD[157] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[158] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[159] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[160] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[161] = 32'b101000_00000000000000000001011010; // jal mod
	HD[162] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[163] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[164] = 32'b000011_00010_00010_0000000000110000; // addi 2 2 48
	HD[165] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[166] = 32'b001011_00000000000000000010101001; // jump _IfExit5_
	HD[167] = 32'b000101_00000_00010_0000000000100000; // li 2 32 / _ElseBegin5_
	HD[168] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[169] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _IfExit5_
	HD[170] = 32'b000101_00000_00011_0000000000010000; // li 3 16
	HD[171] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[172] = 32'b000001_10101_00011_0000000000000010; // lw 3 $fp 2
	HD[173] = 32'b000100_00011_00011_0000000000000010; // subi 3 3 2
	HD[174] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[175] = 32'b000001_10101_00011_0000000000000011; // lw 3 $fp 3
	HD[176] = 32'b100111_00010_00011_00011_00000000000; // lcdwrite 2 3 3
	HD[177] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[178] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[179] = 32'b001111_10110_10111_0000000000000000; // push $ra / print_default_msg
	HD[180] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[181] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[182] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[183] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin6_
	HD[184] = 32'b100111_00000_00000_00000_00001000101; // lcdwrite 0 69
	HD[185] = 32'b100111_00001_00000_00000_00001010010; // lcdwrite 1 82
	HD[186] = 32'b100111_00010_00000_00000_00001010010; // lcdwrite 2 82
	HD[187] = 32'b100111_00011_00000_00000_00001001111; // lcdwrite 3 79
	HD[188] = 32'b100111_00100_00000_00000_00000111010; // lcdwrite 4 58
	HD[189] = 32'b100111_00101_00000_00000_00000100000; // lcdwrite 5 32
	HD[190] = 32'b100111_00110_00000_00000_00001000010; // lcdwrite 6 66
	HD[191] = 32'b100111_00111_00000_00000_00001000001; // lcdwrite 7 65
	HD[192] = 32'b100111_01000_00000_00000_00001000100; // lcdwrite 8 68
	HD[193] = 32'b100111_01001_00000_00000_00000100000; // lcdwrite 9 32
	HD[194] = 32'b100111_01010_00000_00000_00001010110; // lcdwrite 10 86
	HD[195] = 32'b100111_01011_00000_00000_00001000001; // lcdwrite 11 65
	HD[196] = 32'b100111_01100_00000_00000_00001001100; // lcdwrite 12 76
	HD[197] = 32'b100111_01101_00000_00000_00001010101; // lcdwrite 13 85
	HD[198] = 32'b100111_01110_00000_00000_00001000101; // lcdwrite 14 69
	HD[199] = 32'b100111_01111_00000_00000_00000100001; // lcdwrite 15 33
	HD[200] = 32'b001011_00000000000000000101110000; // jump _IfExit6_
	HD[201] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin6_
	HD[202] = 32'b000101_00000_00011_0000000000000010; // li 3 2
	HD[203] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[204] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin7_
	HD[205] = 32'b100111_00000_00000_00000_00001010011; // lcdwrite 0 83
	HD[206] = 32'b100111_00001_00000_00000_00001100101; // lcdwrite 1 101
	HD[207] = 32'b100111_00010_00000_00000_00001101100; // lcdwrite 2 108
	HD[208] = 32'b100111_00011_00000_00000_00001100101; // lcdwrite 3 101
	HD[209] = 32'b100111_00100_00000_00000_00001100011; // lcdwrite 4 99
	HD[210] = 32'b100111_00101_00000_00000_00001101001; // lcdwrite 5 105
	HD[211] = 32'b100111_00110_00000_00000_00001101111; // lcdwrite 6 111
	HD[212] = 32'b100111_00111_00000_00000_00001101110; // lcdwrite 7 110
	HD[213] = 32'b100111_01000_00000_00000_00001100101; // lcdwrite 8 101
	HD[214] = 32'b100111_01001_00000_00000_00000100000; // lcdwrite 9 32
	HD[215] = 32'b100111_01010_00000_00000_00001101111; // lcdwrite 10 111
	HD[216] = 32'b100111_01011_00000_00000_00000100000; // lcdwrite 11 32
	HD[217] = 32'b100111_01100_00000_00000_00001110000; // lcdwrite 12 112
	HD[218] = 32'b100111_01101_00000_00000_00001110010; // lcdwrite 13 114
	HD[219] = 32'b100111_01110_00000_00000_00001101111; // lcdwrite 14 111
	HD[220] = 32'b100111_01111_00000_00000_00001100111; // lcdwrite 15 103
	HD[221] = 32'b001011_00000000000000000101110000; // jump _IfExit7_
	HD[222] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin7_
	HD[223] = 32'b000101_00000_00011_0000000000000011; // li 3 3
	HD[224] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[225] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin8_
	HD[226] = 32'b100111_00000_00000_00000_00001000101; // lcdwrite 0 69
	HD[227] = 32'b100111_00001_00000_00000_00001110010; // lcdwrite 1 114
	HD[228] = 32'b100111_00010_00000_00000_00001110010; // lcdwrite 2 114
	HD[229] = 32'b100111_00011_00000_00000_00001101111; // lcdwrite 3 111
	HD[230] = 32'b100111_00100_00000_00000_00000111010; // lcdwrite 4 58
	HD[231] = 32'b100111_00101_00000_00000_00000100000; // lcdwrite 5 32
	HD[232] = 32'b100111_00110_00000_00000_00001010000; // lcdwrite 6 80
	HD[233] = 32'b100111_00111_00000_00000_00001110010; // lcdwrite 7 114
	HD[234] = 32'b100111_01000_00000_00000_00001101111; // lcdwrite 8 111
	HD[235] = 32'b100111_01001_00000_00000_00001100111; // lcdwrite 9 103
	HD[236] = 32'b100111_01010_00000_00000_00000101110; // lcdwrite 10 46
	HD[237] = 32'b100111_01011_00000_00000_00000100000; // lcdwrite 11 32
	HD[238] = 32'b100111_01100_00000_00000_00000100000; // lcdwrite 12 32
	HD[239] = 32'b100111_01101_00000_00000_00000100000; // lcdwrite 13 32
	HD[240] = 32'b100111_01110_00000_00000_00000100000; // lcdwrite 14 32
	HD[241] = 32'b100111_01111_00000_00000_00000100000; // lcdwrite 15 32
	HD[242] = 32'b001011_00000000000000000101110000; // jump _IfExit8_
	HD[243] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin8_
	HD[244] = 32'b000101_00000_00011_0000000000000100; // li 3 4
	HD[245] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[246] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin9_
	HD[247] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[248] = 32'b100111_10001_00000_00000_00001101110; // lcdwrite 17 110
	HD[249] = 32'b100111_10010_00000_00000_00001100001; // lcdwrite 18 97
	HD[250] = 32'b100111_10011_00000_00000_00001101111; // lcdwrite 19 111
	HD[251] = 32'b100111_10100_00000_00000_00000100000; // lcdwrite 20 32
	HD[252] = 32'b100111_10101_00000_00000_00001100101; // lcdwrite 21 101
	HD[253] = 32'b100111_10110_00000_00000_00001101110; // lcdwrite 22 110
	HD[254] = 32'b100111_10111_00000_00000_00001100011; // lcdwrite 23 99
	HD[255] = 32'b100111_11000_00000_00000_00001101111; // lcdwrite 24 111
	HD[256] = 32'b100111_11001_00000_00000_00001101110; // lcdwrite 25 110
	HD[257] = 32'b100111_11010_00000_00000_00001110100; // lcdwrite 26 116
	HD[258] = 32'b100111_11011_00000_00000_00001110010; // lcdwrite 27 114
	HD[259] = 32'b100111_11100_00000_00000_00001100001; // lcdwrite 28 97
	HD[260] = 32'b100111_11101_00000_00000_00001100100; // lcdwrite 29 100
	HD[261] = 32'b100111_11110_00000_00000_00001101111; // lcdwrite 30 111
	HD[262] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[263] = 32'b001011_00000000000000000101110000; // jump _IfExit9_
	HD[264] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin9_
	HD[265] = 32'b000101_00000_00011_0000000000000101; // li 3 5
	HD[266] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[267] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin10_
	HD[268] = 32'b100111_00000_00000_00000_00000100000; // lcdwrite 0 32
	HD[269] = 32'b100111_00001_00000_00000_00001010000; // lcdwrite 1 80
	HD[270] = 32'b100111_00010_00000_00000_00001110010; // lcdwrite 2 114
	HD[271] = 32'b100111_00011_00000_00000_00001101111; // lcdwrite 3 111
	HD[272] = 32'b100111_00100_00000_00000_00001100111; // lcdwrite 4 103
	HD[273] = 32'b100111_00101_00000_00000_00001110010; // lcdwrite 5 114
	HD[274] = 32'b100111_00110_00000_00000_00001100001; // lcdwrite 6 97
	HD[275] = 32'b100111_00111_00000_00000_00001101101; // lcdwrite 7 109
	HD[276] = 32'b100111_01000_00000_00000_00001100001; // lcdwrite 8 97
	HD[277] = 32'b100111_01001_00000_00000_00000100000; // lcdwrite 9 32
	HD[278] = 32'b100111_01010_00000_00000_00000100000; // lcdwrite 10 32
	HD[279] = 32'b100111_01011_00000_00000_00000100000; // lcdwrite 11 32
	HD[280] = 32'b100111_01100_00000_00000_00000100000; // lcdwrite 12 32
	HD[281] = 32'b100111_01101_00000_00000_00000100000; // lcdwrite 13 32
	HD[282] = 32'b100111_01110_00000_00000_00000100000; // lcdwrite 14 32
	HD[283] = 32'b100111_01111_00000_00000_00000100000; // lcdwrite 15 32
	HD[284] = 32'b001011_00000000000000000101110000; // jump _IfExit10_
	HD[285] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin10_
	HD[286] = 32'b000101_00000_00011_0000000000000110; // li 3 6
	HD[287] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[288] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin11_
	HD[289] = 32'b100111_10000_00000_00000_00001001001; // lcdwrite 16 73
	HD[290] = 32'b100111_10001_00000_00000_00001000100; // lcdwrite 17 68
	HD[291] = 32'b100111_10010_00000_00000_00000100000; // lcdwrite 18 32
	HD[292] = 32'b100111_10011_00000_00000_00001100100; // lcdwrite 19 100
	HD[293] = 32'b100111_10100_00000_00000_00001100101; // lcdwrite 20 101
	HD[294] = 32'b100111_10101_00000_00000_00001110110; // lcdwrite 21 118
	HD[295] = 32'b100111_10110_00000_00000_00001100101; // lcdwrite 22 101
	HD[296] = 32'b100111_10111_00000_00000_00000100000; // lcdwrite 23 32
	HD[297] = 32'b100111_11000_00000_00000_00001110011; // lcdwrite 24 115
	HD[298] = 32'b100111_11001_00000_00000_00001100101; // lcdwrite 25 101
	HD[299] = 32'b100111_11010_00000_00000_00001110010; // lcdwrite 26 114
	HD[300] = 32'b100111_11011_00000_00000_00000100000; // lcdwrite 27 32
	HD[301] = 32'b100111_11100_00000_00000_00000111110; // lcdwrite 28 62
	HD[302] = 32'b100111_11101_00000_00000_00000100000; // lcdwrite 29 32
	HD[303] = 32'b100111_11110_00000_00000_00000110000; // lcdwrite 30 48
	HD[304] = 32'b100111_11111_00000_00000_00000100001; // lcdwrite 31 33
	HD[305] = 32'b001011_00000000000000000101110000; // jump _IfExit11_
	HD[306] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin11_
	HD[307] = 32'b000101_00000_00011_0000000000000111; // li 3 7
	HD[308] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[309] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin12_
	HD[310] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[311] = 32'b100111_10001_00000_00000_00001101010; // lcdwrite 17 106
	HD[312] = 32'b100111_10010_00000_00000_00001100001; // lcdwrite 18 97
	HD[313] = 32'b100111_10011_00000_00000_00000100000; // lcdwrite 19 32
	HD[314] = 32'b100111_10100_00000_00000_00001110101; // lcdwrite 20 117
	HD[315] = 32'b100111_10101_00000_00000_00001110011; // lcdwrite 21 115
	HD[316] = 32'b100111_10110_00000_00000_00001100001; // lcdwrite 22 97
	HD[317] = 32'b100111_10111_00000_00000_00000100000; // lcdwrite 23 32
	HD[318] = 32'b100111_11000_00000_00000_00001100101; // lcdwrite 24 101
	HD[319] = 32'b100111_11001_00000_00000_00001110011; // lcdwrite 25 115
	HD[320] = 32'b100111_11010_00000_00000_00001110011; // lcdwrite 26 115
	HD[321] = 32'b100111_11011_00000_00000_00001100101; // lcdwrite 27 101
	HD[322] = 32'b100111_11100_00000_00000_00000100000; // lcdwrite 28 32
	HD[323] = 32'b100111_11101_00000_00000_00001001001; // lcdwrite 29 73
	HD[324] = 32'b100111_11110_00000_00000_00001000100; // lcdwrite 30 68
	HD[325] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[326] = 32'b001011_00000000000000000101110000; // jump _IfExit12_
	HD[327] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin12_
	HD[328] = 32'b000101_00000_00011_0000000000001000; // li 3 8
	HD[329] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[330] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin13_
	HD[331] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[332] = 32'b100111_10001_00000_00000_00001110011; // lcdwrite 17 115
	HD[333] = 32'b100111_10010_00000_00000_00001100101; // lcdwrite 18 101
	HD[334] = 32'b100111_10011_00000_00000_00001101110; // lcdwrite 19 110
	HD[335] = 32'b100111_10100_00000_00000_00001100100; // lcdwrite 20 100
	HD[336] = 32'b100111_10101_00000_00000_00001101111; // lcdwrite 21 111
	HD[337] = 32'b100111_10110_00000_00000_00000100000; // lcdwrite 22 32
	HD[338] = 32'b100111_10111_00000_00000_00001100101; // lcdwrite 23 101
	HD[339] = 32'b100111_11000_00000_00000_00001111000; // lcdwrite 24 120
	HD[340] = 32'b100111_11001_00000_00000_00001100101; // lcdwrite 25 101
	HD[341] = 32'b100111_11010_00000_00000_00001100011; // lcdwrite 26 99
	HD[342] = 32'b100111_11011_00000_00000_00001110101; // lcdwrite 27 117
	HD[343] = 32'b100111_11100_00000_00000_00001110100; // lcdwrite 28 116
	HD[344] = 32'b100111_11101_00000_00000_00001100001; // lcdwrite 29 97
	HD[345] = 32'b100111_11110_00000_00000_00001100100; // lcdwrite 30 100
	HD[346] = 32'b100111_11111_00000_00000_00001101111; // lcdwrite 31 111
	HD[347] = 32'b001011_00000000000000000101110000; // jump _IfExit13_
	HD[348] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin13_
	HD[349] = 32'b000101_00000_00011_0000000000001001; // li 3 9
	HD[350] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[351] = 32'b000111_00010_00000_0000000000010001; // beq 2 $zero _IfExit14_
	HD[352] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[353] = 32'b100111_10001_00000_00000_00001100110; // lcdwrite 17 102
	HD[354] = 32'b100111_10010_00000_00000_00001101111; // lcdwrite 18 111
	HD[355] = 32'b100111_10011_00000_00000_00001101001; // lcdwrite 19 105
	HD[356] = 32'b100111_10100_00000_00000_00000100000; // lcdwrite 20 32
	HD[357] = 32'b100111_10101_00000_00000_00001100110; // lcdwrite 21 102
	HD[358] = 32'b100111_10110_00000_00000_00001101001; // lcdwrite 22 105
	HD[359] = 32'b100111_10111_00000_00000_00001101110; // lcdwrite 23 110
	HD[360] = 32'b100111_11000_00000_00000_00001100001; // lcdwrite 24 97
	HD[361] = 32'b100111_11001_00000_00000_00001101100; // lcdwrite 25 108
	HD[362] = 32'b100111_11010_00000_00000_00001101001; // lcdwrite 26 105
	HD[363] = 32'b100111_11011_00000_00000_00001111010; // lcdwrite 27 122
	HD[364] = 32'b100111_11100_00000_00000_00001100001; // lcdwrite 28 97
	HD[365] = 32'b100111_11101_00000_00000_00001100100; // lcdwrite 29 100
	HD[366] = 32'b100111_11110_00000_00000_00001101111; // lcdwrite 30 111
	HD[367] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[368] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _IfExit14_ _IfExit13_ _IfExit12_ _IfExit11_ _IfExit10_ _IfExit9_ _IfExit8_ _IfExit7_ _IfExit6_
	HD[369] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[370] = 32'b001111_10110_10111_0000000000000000; // push $ra / load_registradores
	HD[371] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[372] = 32'b000001_00000_00011_0000000000000010; // lw 3 $global 2
	HD[373] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[374] = 32'b000001_00000_00011_0000000000000011; // lw 3 $global 3
	HD[375] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[376] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[377] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[378] = 32'b000001_00010_01010_0000000000001010; // lw 10 2 10
	HD[379] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[380] = 32'b000001_00010_01011_0000000000001011; // lw 11 2 11
	HD[381] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[382] = 32'b000001_00010_01100_0000000000001100; // lw 12 2 12
	HD[383] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[384] = 32'b000001_00010_01101_0000000000001101; // lw 13 2 13
	HD[385] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[386] = 32'b000001_00010_01110_0000000000001110; // lw 14 2 14
	HD[387] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[388] = 32'b000001_00010_01111_0000000000001111; // lw 15 2 15
	HD[389] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[390] = 32'b000001_00010_10000_0000000000010000; // lw 16 2 16
	HD[391] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[392] = 32'b000001_00010_10001_0000000000010001; // lw 17 2 17
	HD[393] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[394] = 32'b000001_00010_10010_0000000000010010; // lw 18 2 18
	HD[395] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[396] = 32'b000001_00010_10011_0000000000010011; // lw 19 2 19
	HD[397] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[398] = 32'b000001_00010_11001_0000000000011001; // lw 25 2 25
	HD[399] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[400] = 32'b000001_00010_11010_0000000000011010; // lw 26 2 26
	HD[401] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[402] = 32'b000001_00010_11011_0000000000011011; // lw 27 2 27
	HD[403] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[404] = 32'b000001_00010_11100_0000000000011100; // lw 28 2 28
	HD[405] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[406] = 32'b000001_00010_11101_0000000000011101; // lw 29 2 29
	HD[407] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[408] = 32'b000001_00010_11110_0000000000011110; // lw 30 2 30
	HD[409] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[410] = 32'b000001_00010_11111_0000000000011111; // lw 31 2 31
	HD[411] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[412] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[413] = 32'b001111_10110_10111_0000000000000000; // push $ra / store_registradores
	HD[414] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[415] = 32'b000001_00000_00011_0000000000000010; // lw 3 $global 2
	HD[416] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[417] = 32'b000001_00000_00011_0000000000000011; // lw 3 $global 3
	HD[418] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[419] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[420] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[421] = 32'b000010_00010_01010_0000000000001010; // sw 10 2 10
	HD[422] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[423] = 32'b000010_00010_01011_0000000000001011; // sw 11 2 11
	HD[424] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[425] = 32'b000010_00010_01100_0000000000001100; // sw 12 2 12
	HD[426] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[427] = 32'b000010_00010_01101_0000000000001101; // sw 13 2 13
	HD[428] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[429] = 32'b000010_00010_01110_0000000000001110; // sw 14 2 14
	HD[430] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[431] = 32'b000010_00010_01111_0000000000001111; // sw 15 2 15
	HD[432] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[433] = 32'b000010_00010_10000_0000000000010000; // sw 16 2 16
	HD[434] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[435] = 32'b000010_00010_10001_0000000000010001; // sw 17 2 17
	HD[436] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[437] = 32'b000010_00010_10010_0000000000010010; // sw 18 2 18
	HD[438] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[439] = 32'b000010_00010_10011_0000000000010011; // sw 19 2 19
	HD[440] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[441] = 32'b000010_00010_11001_0000000000011001; // sw 25 2 25
	HD[442] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[443] = 32'b000010_00010_11010_0000000000011010; // sw 26 2 26
	HD[444] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[445] = 32'b000010_00010_11011_0000000000011011; // sw 27 2 27
	HD[446] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[447] = 32'b000010_00010_11100_0000000000011100; // sw 28 2 28
	HD[448] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[449] = 32'b000010_00010_11101_0000000000011101; // sw 29 2 29
	HD[450] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[451] = 32'b000010_00010_11110_0000000000011110; // sw 30 2 30
	HD[452] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[453] = 32'b000010_00010_11111_0000000000011111; // sw 31 2 31
	HD[454] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[455] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[456] = 32'b001111_10110_10111_0000000000000000; // push $ra / organiza_fila_pronto
	HD[457] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[458] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[459] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
	HD[460] = 32'b000111_00010_00000_0000000000011010; // beq 2 $zero _IfExit15_
	HD[461] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin2_
	HD[462] = 32'b000001_00000_00011_0000000000001000; // lw 3 $global 8
	HD[463] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[464] = 32'b000111_00010_00000_0000000000001100; // beq 2 $zero _WhileExit2_
	HD[465] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[466] = 32'b000000_00010_00000_00010_00000_000101; // add 2 2 $global
	HD[467] = 32'b000001_00010_00010_0000000000001001; // lw 2 2 9
	HD[468] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[469] = 32'b000100_00011_00011_0000000000000001; // subi 3 3 1
	HD[470] = 32'b000000_00011_00000_00011_00000_000101; // add 3 3 $global
	HD[471] = 32'b000010_00011_00010_0000000000001001; // sw 2 3 9
	HD[472] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[473] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[474] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[475] = 32'b001011_00000000000000000111001101; // jump _WhileBegin2_
	HD[476] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileExit2_
	HD[477] = 32'b000001_00000_00011_0000000000000111; // lw 3 $global 7
	HD[478] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
	HD[479] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[480] = 32'b000111_00010_00000_0000000000000110; // beq 2 $zero _IfExit16_
	HD[481] = 32'b000001_00000_00010_0000000000010100; // lw 2 $global 20
	HD[482] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[483] = 32'b000100_00011_00011_0000000000000001; // subi 3 3 1
	HD[484] = 32'b000000_00011_00000_00011_00000_000101; // add 3 3 $global
	HD[485] = 32'b000010_00011_00010_0000000000001001; // sw 2 3 9
	HD[486] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _IfExit16_ _IfExit15_
	HD[487] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[488] = 32'b001111_10110_10111_0000000000000000; // push $ra / fila_existe_processo
	HD[489] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[490] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[491] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _WhileBegin3_
	HD[492] = 32'b000001_00000_00011_0000000000001000; // lw 3 $global 8
	HD[493] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[494] = 32'b000111_00010_00000_0000000000001111; // beq 2 $zero _WhileExit3_
	HD[495] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[496] = 32'b000000_00010_00000_00010_00000_000101; // add 2 2 $global
	HD[497] = 32'b000001_00010_00010_0000000000001001; // lw 2 2 9
	HD[498] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[499] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[500] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _IfExit17_
	HD[501] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[502] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[503] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[504] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[505] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _IfExit17_
	HD[506] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[507] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[508] = 32'b001011_00000000000000000111101011; // jump _WhileBegin3_
	HD[509] = 32'b000001_00000_00010_0000000000010110; // lw 2 $global 22 / _WhileExit3_
	HD[510] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[511] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[512] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[513] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[514] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[515] = 32'b001111_10110_10111_0000000000000000; // push $ra / remove_processo_fila_pronto
	HD[516] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[517] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[518] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _WhileBegin4_
	HD[519] = 32'b000001_00000_00011_0000000000001000; // lw 3 $global 8
	HD[520] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[521] = 32'b000111_00010_00000_0000000000010100; // beq 2 $zero _WhileExit4_
	HD[522] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[523] = 32'b000000_00010_00000_00010_00000_000101; // add 2 2 $global
	HD[524] = 32'b000001_00010_00010_0000000000001001; // lw 2 2 9
	HD[525] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[526] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[527] = 32'b000111_00010_00000_0000000000001010; // beq 2 $zero _IfExit18_
	HD[528] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[529] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[530] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[531] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[532] = 32'b101000_00000000000000000111001000; // jal organiza_fila_pronto
	HD[533] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[534] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8
	HD[535] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[536] = 32'b000010_00000_00010_0000000000001000; // sw 2 $global 8
	HD[537] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _IfExit18_
	HD[538] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[539] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[540] = 32'b001011_00000000000000001000000110; // jump _WhileBegin4_
	HD[541] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _WhileExit4_
	HD[542] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[543] = 32'b001111_10110_10111_0000000000000000; // push $ra / insere_processo_fila_pronto
	HD[544] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[545] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[546] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8
	HD[547] = 32'b000001_00000_00011_0000000000000111; // lw 3 $global 7
	HD[548] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[549] = 32'b000111_00010_00000_0000000000010001; // beq 2 $zero _IfExit19_
	HD[550] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[551] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[552] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[553] = 32'b101000_00000000000000000111101000; // jal fila_existe_processo
	HD[554] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[555] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[556] = 32'b000001_00000_00011_0000000000010110; // lw 3 $global 22
	HD[557] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[558] = 32'b000111_00010_00000_0000000000001000; // beq 2 $zero _IfExit20_
	HD[559] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[560] = 32'b000001_00000_00011_0000000000001000; // lw 3 $global 8
	HD[561] = 32'b000000_00011_00000_00011_00000_000101; // add 3 3 $global
	HD[562] = 32'b000010_00011_00010_0000000000001001; // sw 2 3 9
	HD[563] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8
	HD[564] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[565] = 32'b000010_00000_00010_0000000000001000; // sw 2 $global 8
	HD[566] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _IfExit20_ _IfExit19_
	HD[567] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[568] = 32'b001111_10110_10111_0000000000000000; // push $ra / fila_proximo
	HD[569] = 32'b000001_00000_00010_0000000000001001; // lw 2 $global 9
	HD[570] = 32'b000001_00000_00011_0000000000010100; // lw 3 $global 20
	HD[571] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[572] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[573] = 32'b000111_00010_00000_0000000000001111; // beq 2 $zero _IfExit21_
	HD[574] = 32'b000001_00000_00010_0000000000001001; // lw 2 $global 9
	HD[575] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[576] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[577] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[578] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[579] = 32'b101000_00000000000000000111001000; // jal organiza_fila_pronto
	HD[580] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[581] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8
	HD[582] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[583] = 32'b000010_00000_00010_0000000000001000; // sw 2 $global 8
	HD[584] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[585] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[586] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[587] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[588] = 32'b000001_00000_00010_0000000000010101; // lw 2 $global 21 / _IfExit21_
	HD[589] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[590] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[591] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[592] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[593] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[594] = 32'b001111_10110_10111_0000000000000000; // push $ra / fila_passa_vez
	HD[595] = 32'b000001_00000_00010_0000000000001001; // lw 2 $global 9
	HD[596] = 32'b000001_00000_00011_0000000000010100; // lw 3 $global 20
	HD[597] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[598] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[599] = 32'b000111_00010_00000_0000000000001101; // beq 2 $zero _IfExit22_
	HD[600] = 32'b000001_00000_00010_0000000000001001; // lw 2 $global 9
	HD[601] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[602] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[603] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[604] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[605] = 32'b101000_00000000000000000111001000; // jal organiza_fila_pronto
	HD[606] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[607] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[608] = 32'b000001_00000_00011_0000000000001000; // lw 3 $global 8
	HD[609] = 32'b000100_00011_00011_0000000000000001; // subi 3 3 1
	HD[610] = 32'b000000_00011_00000_00011_00000_000101; // add 3 3 $global
	HD[611] = 32'b000010_00011_00010_0000000000001001; // sw 2 3 9
	HD[612] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _IfExit22_
	HD[613] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[614] = 32'b001111_10110_10111_0000000000000000; // push $ra / posicao_programa
	HD[615] = 32'b000001_00000_00010_0000000000010111; // lw 2 $global 23
	HD[616] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[617] = 32'b000001_00000_00010_0000000000011110; // lw 2 $global 30
	HD[618] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[619] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[620] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[621] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _WhileBegin5_
	HD[622] = 32'b000001_00000_00011_0000000000000000; // lw 3 $global 0
	HD[623] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[624] = 32'b000111_00010_00000_0000000000011100; // beq 2 $zero _WhileExit5_
	HD[625] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[626] = 32'b000001_10101_00011_0000000000000001; // lw 3 $fp 1
	HD[627] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[628] = 32'b000010_10101_00010_0000000000000101; // sw 2 $fp 5
	HD[629] = 32'b000001_10101_00010_0000000000000101; // lw 2 $fp 5
	HD[630] = 32'b000001_00000_00011_0000000000011101; // lw 3 $global 29
	HD[631] = 32'b100100_00010_00011_00010_00000_000000; // hdtoreg 2 2 3
	HD[632] = 32'b000001_00000_00011_0000000000011000; // lw 3 $global 24
	HD[633] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[634] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[635] = 32'b000111_00010_00000_0000000000001101; // beq 2 $zero _IfExit23_
	HD[636] = 32'b000001_10101_00010_0000000000000101; // lw 2 $fp 5
	HD[637] = 32'b000001_10101_00011_0000000000000011; // lw 3 $fp 3
	HD[638] = 32'b100100_00010_00011_00010_00000_000000; // hdtoreg 2 2 3
	HD[639] = 32'b000010_10101_00010_0000000000000100; // sw 2 $fp 4
	HD[640] = 32'b000001_10101_00010_0000000000000100; // lw 2 $fp 4
	HD[641] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[642] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[643] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _IfExit24_
	HD[644] = 32'b000001_10101_00010_0000000000000101; // lw 2 $fp 5
	HD[645] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[646] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[647] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[648] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _IfExit24_ _IfExit23_
	HD[649] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[650] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[651] = 32'b001011_00000000000000001001101101; // jump _WhileBegin5_
	HD[652] = 32'b000001_00000_00010_0000000000011001; // lw 2 $global 25 / _WhileExit5_
	HD[653] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[654] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[655] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[656] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[657] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[658] = 32'b001111_10110_10111_0000000000000000; // push $ra / posicao_livre_programa
	HD[659] = 32'b000001_00000_00010_0000000000010111; // lw 2 $global 23
	HD[660] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[661] = 32'b000001_00000_00010_0000000000011101; // lw 2 $global 29
	HD[662] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[663] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[664] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[665] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin6_
	HD[666] = 32'b000001_00000_00011_0000000000000000; // lw 3 $global 0
	HD[667] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[668] = 32'b000111_00010_00000_0000000000010011; // beq 2 $zero _WhileExit6_
	HD[669] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[670] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[671] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[672] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[673] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3
	HD[674] = 32'b000001_10101_00011_0000000000000010; // lw 3 $fp 2
	HD[675] = 32'b100100_00010_00011_00010_00000_000000; // hdtoreg 2 2 3
	HD[676] = 32'b000001_00000_00011_0000000000011000; // lw 3 $global 24
	HD[677] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[678] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _IfExit25_
	HD[679] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3
	HD[680] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[681] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[682] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[683] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _IfExit25_
	HD[684] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[685] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[686] = 32'b001011_00000000000000001010011001; // jump _WhileBegin6_
	HD[687] = 32'b000001_00000_00010_0000000000011010; // lw 2 $global 26 / _WhileExit6_
	HD[688] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[689] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[690] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[691] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[692] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[693] = 32'b001111_10110_10111_0000000000000000; // push $ra / tamanho_programa
	HD[694] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[695] = 32'b000011_10101_10101_0000000000000011; // addi $fp $fp 3
	HD[696] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[697] = 32'b101000_00000000000000001001100110; // jal posicao_programa
	HD[698] = 32'b000100_10101_10101_0000000000000011; // subi $fp $fp 3
	HD[699] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[700] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[701] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[702] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[703] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[704] = 32'b000111_00010_00000_0000000000000110; // beq 2 $zero _IfExit26_
	HD[705] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[706] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[707] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[708] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[709] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[710] = 32'b000001_00000_00010_0000000000100000; // lw 2 $global 32 / _IfExit26_
	HD[711] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[712] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[713] = 32'b000001_00000_00011_0000000000011111; // lw 3 $global 31
	HD[714] = 32'b100100_00010_00011_00010_00000_000000; // hdtoreg 2 2 3
	HD[715] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[716] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[717] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[718] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[719] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[720] = 32'b001111_10110_10111_0000000000000000; // push $ra / carrega_programa_memoria_inst
	HD[721] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[722] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[723] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[724] = 32'b000011_10101_10101_0000000000000101; // addi $fp $fp 5
	HD[725] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[726] = 32'b101000_00000000000000001001100110; // jal posicao_programa
	HD[727] = 32'b000100_10101_10101_0000000000000101; // subi $fp $fp 5
	HD[728] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[729] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[730] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[731] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[732] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[733] = 32'b000111_00010_00000_0000000000000110; // beq 2 $zero _IfExit27_
	HD[734] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[735] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[736] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[737] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[738] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[739] = 32'b000001_00000_00010_0000000000100000; // lw 2 $global 32 / _IfExit27_
	HD[740] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[741] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[742] = 32'b000001_00000_00011_0000000000011111; // lw 3 $global 31
	HD[743] = 32'b100100_00010_00011_00010_00000_000000; // hdtoreg 2 2 3
	HD[744] = 32'b000010_10101_00010_0000000000000100; // sw 2 $fp 4
	HD[745] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _WhileBegin7_
	HD[746] = 32'b000001_10101_00011_0000000000000100; // lw 3 $fp 4
	HD[747] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[748] = 32'b000111_00010_00000_0000000000001101; // beq 2 $zero _WhileExit7_
	HD[749] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[750] = 32'b000001_10101_00011_0000000000000011; // lw 3 $fp 3
	HD[751] = 32'b000001_10101_00100_0000000000000001; // lw 4 $fp 1
	HD[752] = 32'b000000_00011_00100_00011_00000_000101; // add 3 3 4
	HD[753] = 32'b000001_00000_00100_0000000000000001; // lw 4 $global 1
	HD[754] = 32'b000001_10101_00101_0000000000000001; // lw 5 $fp 1
	HD[755] = 32'b000000_00100_00101_00100_00000_000101; // add 4 4 5
	HD[756] = 32'b100011_00010_00011_00100_00000_000000; // hdtoinst 4 2 3
	HD[757] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[758] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[759] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[760] = 32'b001011_00000000000000001011101001; // jump _WhileBegin7_
	HD[761] = 32'b000001_10101_00010_0000000000000100; // lw 2 $fp 4 / _WhileExit7_
	HD[762] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[763] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[764] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[765] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[766] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[767] = 32'b001111_10110_10111_0000000000000000; // push $ra / cria_programa
	HD[768] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[769] = 32'b000011_10101_10101_0000000000000111; // addi $fp $fp 7
	HD[770] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[771] = 32'b101000_00000000000000001001100110; // jal posicao_programa
	HD[772] = 32'b000100_10101_10101_0000000000000111; // subi $fp $fp 7
	HD[773] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[774] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[775] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[776] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[777] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[778] = 32'b000111_00010_00000_0000000000111101; // beq 2 $zero _IfExit28_
	HD[779] = 32'b000011_10101_10101_0000000000000111; // addi $fp $fp 7
	HD[780] = 32'b101000_00000000000000001010010010; // jal posicao_livre_programa
	HD[781] = 32'b000100_10101_10101_0000000000000111; // subi $fp $fp 7
	HD[782] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[783] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[784] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[785] = 32'b000001_00000_00011_0000000000011101; // lw 3 $global 29
	HD[786] = 32'b000101_00000_00100_0000000000000001; // li 4 1
	HD[787] = 32'b100101_00010_00011_00100_00000_000000; // regtohd 4 2 3
	HD[788] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[789] = 32'b000001_00000_00011_0000000000011110; // lw 3 $global 30
	HD[790] = 32'b000001_10101_00100_0000000000000000; // lw 4 $fp 0
	HD[791] = 32'b100101_00010_00011_00100_00000_000000; // regtohd 4 2 3
	HD[792] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[793] = 32'b000001_00000_00011_0000000000011111; // lw 3 $global 31
	HD[794] = 32'b000001_10101_00100_0000000000000001; // lw 4 $fp 1
	HD[795] = 32'b100101_00010_00011_00100_00000_000000; // regtohd 4 2 3
	HD[796] = 32'b000001_00000_00010_0000000000011100; // lw 2 $global 28
	HD[797] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[798] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[799] = 32'b000001_00000_00011_0000000000011100; // lw 3 $global 28
	HD[800] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[801] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[802] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[803] = 32'b000010_10101_00010_0000000000000110; // sw 2 $fp 6
	HD[804] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3 / _WhileBegin8_
	HD[805] = 32'b000001_10101_00011_0000000000000001; // lw 3 $fp 1
	HD[806] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[807] = 32'b000111_00010_00000_0000000000011101; // beq 2 $zero _WhileExit8_
	HD[808] = 32'b000001_10101_00010_0000000000000110; // lw 2 $fp 6
	HD[809] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[810] = 32'b000101_00000_00100_0000000000001111; // li 4 15
	HD[811] = 32'b000011_10101_10101_0000000000000111; // addi $fp $fp 7
	HD[812] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[813] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[814] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[815] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[816] = 32'b000100_10101_10101_0000000000000111; // subi $fp $fp 7
	HD[817] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[818] = 32'b000010_10101_00010_0000000000000100; // sw 2 $fp 4
	HD[819] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[820] = 32'b000010_10101_00010_0000000000000101; // sw 2 $fp 5
	HD[821] = 32'b000001_10101_00010_0000000000000100; // lw 2 $fp 4
	HD[822] = 32'b000001_10101_00011_0000000000000101; // lw 3 $fp 5
	HD[823] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[824] = 32'b000010_10101_00010_0000000000000100; // sw 2 $fp 4
	HD[825] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[826] = 32'b000001_10101_00011_0000000000000011; // lw 3 $fp 3
	HD[827] = 32'b000001_10101_00100_0000000000000100; // lw 4 $fp 4
	HD[828] = 32'b100101_00010_00011_00100_00000_000000; // regtohd 4 2 3
	HD[829] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3
	HD[830] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[831] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[832] = 32'b000001_10101_00010_0000000000000110; // lw 2 $fp 6
	HD[833] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[834] = 32'b000010_10101_00010_0000000000000110; // sw 2 $fp 6
	HD[835] = 32'b001011_00000000000000001100100100; // jump _WhileBegin8_
	HD[836] = 32'b000101_00000_10100_0000000000000001; // li $rv 1 / _WhileExit8_
	HD[837] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[838] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[839] = 32'b000001_00000_00010_0000000000011011; // lw 2 $global 27 / _IfExit28_
	HD[840] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[841] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[842] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[843] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[844] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[845] = 32'b001111_10110_10111_0000000000000000; // push $ra / deleta_programa
	HD[846] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[847] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[848] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[849] = 32'b101000_00000000000000001001100110; // jal posicao_programa
	HD[850] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[851] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[852] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[853] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[854] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[855] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[856] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[857] = 32'b000111_00010_00000_0000000000001000; // beq 2 $zero _IfExit29_
	HD[858] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[859] = 32'b000001_00000_00011_0000000000011101; // lw 3 $global 29
	HD[860] = 32'b000101_00000_00100_0000000000000000; // li 4 0
	HD[861] = 32'b100101_00010_00011_00100_00000_000000; // regtohd 4 2 3
	HD[862] = 32'b000101_00000_10100_0000000000000001; // li $rv 1
	HD[863] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[864] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[865] = 32'b000001_00000_00010_0000000000011001; // lw 2 $global 25 / _IfExit29_
	HD[866] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[867] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[868] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[869] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[870] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[871] = 32'b001111_10110_10111_0000000000000000; // push $ra / renomear_programa
	HD[872] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[873] = 32'b000011_10101_10101_0000000000000011; // addi $fp $fp 3
	HD[874] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[875] = 32'b101000_00000000000000001001100110; // jal posicao_programa
	HD[876] = 32'b000100_10101_10101_0000000000000011; // subi $fp $fp 3
	HD[877] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[878] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[879] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[880] = 32'b000111_00010_00000_0000000000011010; // beq 2 $zero _ElseBegin30_
	HD[881] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[882] = 32'b000011_10101_10101_0000000000000011; // addi $fp $fp 3
	HD[883] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[884] = 32'b101000_00000000000000001001100110; // jal posicao_programa
	HD[885] = 32'b000100_10101_10101_0000000000000011; // subi $fp $fp 3
	HD[886] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[887] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[888] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[889] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[890] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[891] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[892] = 32'b000111_00010_00000_0000000000001001; // beq 2 $zero _ElseBegin31_
	HD[893] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[894] = 32'b000001_00000_00011_0000000000011110; // lw 3 $global 30
	HD[895] = 32'b000001_10101_00100_0000000000000001; // lw 4 $fp 1
	HD[896] = 32'b100101_00010_00011_00100_00000_000000; // regtohd 4 2 3
	HD[897] = 32'b000101_00000_10100_0000000000000001; // li $rv 1
	HD[898] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[899] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[900] = 32'b001011_00000000000000001110001001; // jump _IfExit31_
	HD[901] = 32'b000001_00000_00010_0000000000011001; // lw 2 $global 25 / _ElseBegin31_
	HD[902] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[903] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[904] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[905] = 32'b001011_00000000000000001110001110; // jump _IfExit30_ / _IfExit31_
	HD[906] = 32'b000001_00000_00010_0000000000011011; // lw 2 $global 27 / _ElseBegin30_
	HD[907] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[908] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[909] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[910] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _IfExit30_
	HD[911] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[912] = 32'b001111_10110_10111_0000000000000000; // push $ra / trilha_possui_programa
	HD[913] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[914] = 32'b000001_00000_00011_0000000000010111; // lw 3 $global 23
	HD[915] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[916] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[917] = 32'b000111_00010_00000_0000000000001110; // beq 2 $zero _IfExit32_
	HD[918] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[919] = 32'b000001_00000_00011_0000000000011101; // lw 3 $global 29
	HD[920] = 32'b100100_00010_00011_00010_00000_000000; // hdtoreg 2 2 3
	HD[921] = 32'b000001_00000_00011_0000000000011000; // lw 3 $global 24
	HD[922] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[923] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[924] = 32'b000111_00010_00000_0000000000000111; // beq 2 $zero _IfExit33_
	HD[925] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[926] = 32'b000001_00000_00011_0000000000011110; // lw 3 $global 30
	HD[927] = 32'b100100_00010_00011_00010_00000_000000; // hdtoreg 2 2 3
	HD[928] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[929] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[930] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[931] = 32'b000001_00000_00010_0000000000011001; // lw 2 $global 25 / _IfExit33_ _IfExit32_
	HD[932] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[933] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[934] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[935] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[936] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[937] = 32'b001111_10110_10111_0000000000000000; // push $ra / existe_programa_posicao
	HD[938] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[939] = 32'b000001_00000_00011_0000000000010111; // lw 3 $global 23
	HD[940] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[941] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[942] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[943] = 32'b101000_00000000000000001110010000; // jal trilha_possui_programa
	HD[944] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[945] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[946] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[947] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[948] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[949] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[950] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[951] = 32'b001111_10110_10111_0000000000000000; // push $ra / executa_processos
	HD[952] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[953] = 32'b000010_00000_00010_0000000000000110; // sw 2 $global 6
	HD[954] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8 / _WhileBegin9_
	HD[955] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[956] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
	HD[957] = 32'b000111_00010_00000_0000000001000110; // beq 2 $zero _WhileExit9_
	HD[958] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[959] = 32'b101000_00000000000000001000111000; // jal fila_proximo
	HD[960] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[961] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[962] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[963] = 32'b000101_00000_00010_0000000000000101; // li 2 5
	HD[964] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[965] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[966] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[967] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[968] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[969] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[970] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[971] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[972] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[973] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[974] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[975] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[976] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[977] = 32'b000101_00000_00010_0000000000001000; // li 2 8
	HD[978] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[979] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[980] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[981] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[982] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[983] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[984] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[985] = 32'b101000_00000000000000001011010000; // jal carrega_programa_memoria_inst
	HD[986] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[987] = 32'b000001_00000_00010_0000000000000100; // lw 2 $global 4
	HD[988] = 32'b000001_00000_00011_0000000000000101; // lw 3 $global 5
	HD[989] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[990] = 32'b000000_00010_11110_00000_00000_010000; // move 30 2
	HD[991] = 32'b000001_00000_00010_0000000000000010; // lw 2 $global 2
	HD[992] = 32'b000001_00000_00011_0000000000000011; // lw 3 $global 3
	HD[993] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[994] = 32'b000001_00000_00011_0000000000000101; // lw 3 $global 5
	HD[995] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[996] = 32'b000000_00010_11011_00000_00000_010000; // move 27 2
	HD[997] = 32'b000001_00000_00010_0000000000000001; // lw 2 $global 1
	HD[998] = 32'b000000_00010_00000_00000_00000_010100; // jr 2
	HD[999] = 32'b00000000000000000000000000000000; // noop / _label1_
	HD[1000] = 32'b000101_00000_00010_0000000000000101; // li 2 5
	HD[1001] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[1002] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1003] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1004] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[1005] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[1006] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1007] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[1008] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[1009] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[1010] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1011] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1012] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[1013] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[1014] = 32'b000101_00000_00010_0000000000001001; // li 2 9
	HD[1015] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[1016] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1017] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1018] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[1019] = 32'b000101_00000_00010_0000000000000011; // li 2 3
	HD[1020] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1021] = 32'b000011_10101_10101_0000000000000001; // addi $fp $fp 1
	HD[1022] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1023] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1024] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1025] = 32'b000100_10101_10101_0000000000000001; // subi $fp $fp 1
	HD[1026] = 32'b001011_00000000000000001110111010; // jump _WhileBegin9_
	HD[1027] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _WhileExit9_
	HD[1028] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[1029] = 32'b001111_10110_10111_0000000000000000; // push $ra / executa_processos_preemptivo
	HD[1030] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[1031] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1032] = 32'b000010_10101_00010_0000000000000100; // sw 2 $fp 4
	HD[1033] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin10_
	HD[1034] = 32'b000001_00000_00011_0000000000000111; // lw 3 $global 7
	HD[1035] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[1036] = 32'b000111_00010_00000_0000000000001111; // beq 2 $zero _WhileExit10_
	HD[1037] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[1038] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[1039] = 32'b000000_00011_10101_00011_00000_000101; // add 3 3 $fp
	HD[1040] = 32'b000010_00011_00010_0000000000000101; // sw 2 3 5
	HD[1041] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[1042] = 32'b000000_00010_00000_00010_00000_000101; // add 2 2 $global
	HD[1043] = 32'b000001_00010_00010_0000000000001001; // lw 2 2 9
	HD[1044] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[1045] = 32'b000000_00011_10101_00011_00000_000101; // add 3 3 $fp
	HD[1046] = 32'b000010_00011_00010_0000000000001111; // sw 2 3 15
	HD[1047] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[1048] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[1049] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1050] = 32'b001011_00000000000000010000001001; // jump _WhileBegin10_
	HD[1051] = 32'b000101_00000_00010_0000000000000010; // li 2 2 / _WhileExit10_
	HD[1052] = 32'b000010_00000_00010_0000000000000110; // sw 2 $global 6
	HD[1053] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8 / _WhileBegin11_
	HD[1054] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1055] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
	HD[1056] = 32'b000111_00010_00000_0000000011010011; // beq 2 $zero _WhileExit11_
	HD[1057] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[1058] = 32'b000010_00000_00010_0000000000010011; // sw 2 $global 19
	HD[1059] = 32'b000001_00000_00010_0000000000001001; // lw 2 $global 9
	HD[1060] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[1061] = 32'b100110_00000000000000000000000000; // lcdclean
	HD[1062] = 32'b000001_10101_00010_0000000000000100; // lw 2 $fp 4
	HD[1063] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[1064] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1065] = 32'b000111_00010_00000_0000000000111110; // beq 2 $zero _IfExit34_
	HD[1066] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8
	HD[1067] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[1068] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1069] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[1070] = 32'b000111_00010_00000_0000000000111001; // beq 2 $zero _IfExit35_
	HD[1071] = 32'b100111_00000_00000_00000_00001010010; // lcdwrite 0 82
	HD[1072] = 32'b100111_00001_00000_00000_00001100101; // lcdwrite 1 101
	HD[1073] = 32'b100111_00010_00000_00000_00001100001; // lcdwrite 2 97
	HD[1074] = 32'b100111_00011_00000_00000_00001101100; // lcdwrite 3 108
	HD[1075] = 32'b100111_00100_00000_00000_00001101001; // lcdwrite 4 105
	HD[1076] = 32'b100111_00101_00000_00000_00001111010; // lcdwrite 5 122
	HD[1077] = 32'b100111_00110_00000_00000_00001100001; // lcdwrite 6 97
	HD[1078] = 32'b100111_00111_00000_00000_00001101110; // lcdwrite 7 110
	HD[1079] = 32'b100111_01000_00000_00000_00001100100; // lcdwrite 8 100
	HD[1080] = 32'b100111_01001_00000_00000_00001101111; // lcdwrite 9 111
	HD[1081] = 32'b100111_01011_00000_00000_00001110100; // lcdwrite 11 116
	HD[1082] = 32'b100111_01100_00000_00000_00001110010; // lcdwrite 12 114
	HD[1083] = 32'b100111_01101_00000_00000_00001101111; // lcdwrite 13 111
	HD[1084] = 32'b100111_01110_00000_00000_00001100011; // lcdwrite 14 99
	HD[1085] = 32'b100111_01111_00000_00000_00001100001; // lcdwrite 15 97
	HD[1086] = 32'b100111_10000_00000_00000_00001100100; // lcdwrite 16 100
	HD[1087] = 32'b100111_10001_00000_00000_00001100101; // lcdwrite 17 101
	HD[1088] = 32'b100111_10011_00000_00000_00001000011; // lcdwrite 19 67
	HD[1089] = 32'b100111_10100_00000_00000_00001101111; // lcdwrite 20 111
	HD[1090] = 32'b100111_10101_00000_00000_00001101110; // lcdwrite 21 110
	HD[1091] = 32'b100111_10110_00000_00000_00001110100; // lcdwrite 22 116
	HD[1092] = 32'b100111_10111_00000_00000_00001100101; // lcdwrite 23 101
	HD[1093] = 32'b100111_11000_00000_00000_00001111000; // lcdwrite 24 120
	HD[1094] = 32'b100111_11001_00000_00000_00001110100; // lcdwrite 25 116
	HD[1095] = 32'b100111_11010_00000_00000_00001101111; // lcdwrite 26 111
	HD[1096] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1097] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1098] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1099] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1100] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1101] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1102] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1103] = 32'b100111_11100_00000_00000_00000101110; // lcdwrite 28 46
	HD[1104] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1105] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1106] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1107] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1108] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1109] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1110] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1111] = 32'b100111_11101_00000_00000_00000101110; // lcdwrite 29 46
	HD[1112] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1113] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1114] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1115] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1116] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1117] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1118] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1119] = 32'b100111_11110_00000_00000_00000101110; // lcdwrite 30 46
	HD[1120] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1121] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1122] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1123] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1124] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1125] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1126] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1127] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _IfExit35_ _IfExit34_
	HD[1128] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1129] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1130] = 32'b101000_00000000000000001011010000; // jal carrega_programa_memoria_inst
	HD[1131] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1132] = 32'b000011_10101_00010_0000000000001111; // addi 2 $fp 15
	HD[1133] = 32'b000001_00000_00011_0000000000000111; // lw 3 $global 7
	HD[1134] = 32'b000001_10101_00100_0000000000000001; // lw 4 $fp 1
	HD[1135] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1136] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[1137] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1138] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1139] = 32'b101000_00000000000000000000111101; // jal vetor_existe_valor
	HD[1140] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1141] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[1142] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[1143] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[1144] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3
	HD[1145] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[1146] = 32'b000000_00010_10101_00010_00000_000101; // add 2 2 $fp
	HD[1147] = 32'b000001_00010_00010_0000000000000101; // lw 2 2 5
	HD[1148] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1149] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1150] = 32'b000111_00010_00000_0000000000010111; // beq 2 $zero _ElseBegin36_
	HD[1151] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3
	HD[1152] = 32'b000001_00000_00011_0000000000000100; // lw 3 $global 4
	HD[1153] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[1154] = 32'b000001_00000_00011_0000000000000101; // lw 3 $global 5
	HD[1155] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[1156] = 32'b000000_00010_11110_00000_00000_010000; // move 30 2
	HD[1157] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3
	HD[1158] = 32'b000001_00000_00011_0000000000000010; // lw 3 $global 2
	HD[1159] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[1160] = 32'b000001_00000_00011_0000000000000011; // lw 3 $global 3
	HD[1161] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[1162] = 32'b000001_00000_00011_0000000000000101; // lw 3 $global 5
	HD[1163] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[1164] = 32'b000000_00010_11011_00000_00000_010000; // move 27 2
	HD[1165] = 32'b000001_00000_00010_0000000000000001; // lw 2 $global 1
	HD[1166] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[1167] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1168] = 32'b000001_10101_00011_0000000000000011; // lw 3 $fp 3
	HD[1169] = 32'b000100_00011_00011_0000000000000001; // subi 3 3 1
	HD[1170] = 32'b000000_00011_10101_00011_00000_000101; // add 3 3 $fp
	HD[1171] = 32'b000010_00011_00010_0000000000000101; // sw 2 3 5
	HD[1172] = 32'b001011_00000000000000010010011100; // jump _IfExit36_
	HD[1173] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3 / _ElseBegin36_
	HD[1174] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1175] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1176] = 32'b101000_00000000000000000101110010; // jal load_registradores
	HD[1177] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1178] = 32'b000000_11010_00010_00000_00000_010000; // move 2 26
	HD[1179] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[1180] = 32'b000101_00000_00010_0000000000000101; // li 2 5 / _IfExit36_
	HD[1181] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1182] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1183] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1184] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1185] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[1186] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1187] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[1188] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1189] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[1190] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1191] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1192] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[1193] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1194] = 32'b000101_00000_00010_0000000000001000; // li 2 8
	HD[1195] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1196] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1197] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1198] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1199] = 32'b101010_00000000000000000000000000; // intr_on
	HD[1200] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[1201] = 32'b000000_00010_00000_00000_00000_010100; // jr 2
	HD[1202] = 32'b00000000000000000000000000000000; // noop / _label2_
	HD[1203] = 32'b000001_00000_00010_0000000000010011; // lw 2 $global 19
	HD[1204] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[1205] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1206] = 32'b000111_00010_00000_0000000000010110; // beq 2 $zero _ElseBegin37_
	HD[1207] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1208] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1209] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1210] = 32'b101000_00000000000000000111001000; // jal organiza_fila_pronto
	HD[1211] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1212] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8
	HD[1213] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[1214] = 32'b000010_00000_00010_0000000000001000; // sw 2 $global 8
	HD[1215] = 32'b000101_00000_00010_0000000000001001; // li 2 9
	HD[1216] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1217] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1218] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1219] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1220] = 32'b000101_00000_00010_0000000000000010; // li 2 2
	HD[1221] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1222] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1223] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1224] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1225] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1226] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1227] = 32'b001011_00000000000000010011110000; // jump _IfExit37_
	HD[1228] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3 / _ElseBegin37_
	HD[1229] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1230] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1231] = 32'b101000_00000000000000000110011101; // jal store_registradores
	HD[1232] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1233] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1234] = 32'b101000_00000000000000001001010010; // jal fila_passa_vez
	HD[1235] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1236] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8
	HD[1237] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[1238] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1239] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[1240] = 32'b000111_00010_00000_0000000000011000; // beq 2 $zero _IfExit38_
	HD[1241] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[1242] = 32'b100111_10001_00000_00000_00001100110; // lcdwrite 17 102
	HD[1243] = 32'b100111_10010_00000_00000_00001101111; // lcdwrite 18 111
	HD[1244] = 32'b100111_10011_00000_00000_00001101001; // lcdwrite 19 105
	HD[1245] = 32'b100111_10100_00000_00000_00000100000; // lcdwrite 20 32
	HD[1246] = 32'b100111_10101_00000_00000_00001110000; // lcdwrite 21 112
	HD[1247] = 32'b100111_10110_00000_00000_00001110010; // lcdwrite 22 114
	HD[1248] = 32'b100111_10111_00000_00000_00001100101; // lcdwrite 23 101
	HD[1249] = 32'b100111_11000_00000_00000_00001100101; // lcdwrite 24 101
	HD[1250] = 32'b100111_11001_00000_00000_00001101101; // lcdwrite 25 109
	HD[1251] = 32'b100111_11010_00000_00000_00001110000; // lcdwrite 26 112
	HD[1252] = 32'b100111_11011_00000_00000_00001110100; // lcdwrite 27 116
	HD[1253] = 32'b100111_11100_00000_00000_00001100001; // lcdwrite 28 97
	HD[1254] = 32'b100111_11101_00000_00000_00001100100; // lcdwrite 29 100
	HD[1255] = 32'b100111_11110_00000_00000_00001101111; // lcdwrite 30 111
	HD[1256] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[1257] = 32'b000101_00000_00010_0000000000000010; // li 2 2
	HD[1258] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1259] = 32'b000011_10101_10101_0000000000011001; // addi $fp $fp 25
	HD[1260] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1261] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1262] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1263] = 32'b000100_10101_10101_0000000000011001; // subi $fp $fp 25
	HD[1264] = 32'b000101_00000_00010_0000000000000001; // li 2 1 / _IfExit38_ _IfExit37_
	HD[1265] = 32'b000010_10101_00010_0000000000000100; // sw 2 $fp 4
	HD[1266] = 32'b001011_00000000000000010000011101; // jump _WhileBegin11_
	HD[1267] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _WhileExit11_
	HD[1268] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[1269] = 32'b001111_10110_10111_0000000000000000; // push $ra / seleciona_programas
	HD[1270] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[1271] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[1272] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8
	HD[1273] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1274] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1275] = 32'b000111_00010_00000_0000000100000000; // beq 2 $zero _IfExit39_
	HD[1276] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1277] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1278] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin12_
	HD[1279] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[1280] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1281] = 32'b000111_00010_00000_0000000001101000; // beq 2 $zero _WhileExit12_
	HD[1282] = 32'b100111_00000_00000_00000_00001010011; // lcdwrite 0 83
	HD[1283] = 32'b100111_00001_00000_00000_00001100101; // lcdwrite 1 101
	HD[1284] = 32'b100111_00010_00000_00000_00001101100; // lcdwrite 2 108
	HD[1285] = 32'b100111_00011_00000_00000_00001100101; // lcdwrite 3 101
	HD[1286] = 32'b100111_00100_00000_00000_00001100011; // lcdwrite 4 99
	HD[1287] = 32'b100111_00101_00000_00000_00001101001; // lcdwrite 5 105
	HD[1288] = 32'b100111_00110_00000_00000_00001101111; // lcdwrite 6 111
	HD[1289] = 32'b100111_00111_00000_00000_00001101110; // lcdwrite 7 110
	HD[1290] = 32'b100111_01000_00000_00000_00001100101; // lcdwrite 8 101
	HD[1291] = 32'b100111_01001_00000_00000_00000100000; // lcdwrite 9 32
	HD[1292] = 32'b100111_01010_00000_00000_00001100001; // lcdwrite 10 97
	HD[1293] = 32'b100111_01011_00000_00000_00000100000; // lcdwrite 11 32
	HD[1294] = 32'b100111_01100_00000_00000_00001110001; // lcdwrite 12 113
	HD[1295] = 32'b100111_01101_00000_00000_00001110100; // lcdwrite 13 116
	HD[1296] = 32'b100111_01110_00000_00000_00001100100; // lcdwrite 14 100
	HD[1297] = 32'b100111_01111_00000_00000_00000101110; // lcdwrite 15 46
	HD[1298] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[1299] = 32'b100111_10001_00000_00000_00000100000; // lcdwrite 17 32
	HD[1300] = 32'b100111_10010_00000_00000_00001100100; // lcdwrite 18 100
	HD[1301] = 32'b100111_10011_00000_00000_00001100101; // lcdwrite 19 101
	HD[1302] = 32'b100111_10100_00000_00000_00000100000; // lcdwrite 20 32
	HD[1303] = 32'b100111_10101_00000_00000_00001110000; // lcdwrite 21 112
	HD[1304] = 32'b100111_10110_00000_00000_00001110010; // lcdwrite 22 114
	HD[1305] = 32'b100111_10111_00000_00000_00001101111; // lcdwrite 23 111
	HD[1306] = 32'b100111_11000_00000_00000_00001100111; // lcdwrite 24 103
	HD[1307] = 32'b100111_11001_00000_00000_00001110010; // lcdwrite 25 114
	HD[1308] = 32'b100111_11010_00000_00000_00001100001; // lcdwrite 26 97
	HD[1309] = 32'b100111_11011_00000_00000_00001101101; // lcdwrite 27 109
	HD[1310] = 32'b100111_11100_00000_00000_00001100001; // lcdwrite 28 97
	HD[1311] = 32'b100111_11101_00000_00000_00001110011; // lcdwrite 29 115
	HD[1312] = 32'b100111_11110_00000_00000_00000100000; // lcdwrite 30 32
	HD[1313] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[1314] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[1315] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[1316] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[1317] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1318] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[1319] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[1320] = 32'b000111_00010_00000_0000000000011100; // beq 2 $zero _ElseBegin40_
	HD[1321] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[1322] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[1323] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
	HD[1324] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[1325] = 32'b000111_00010_00000_0000000000000100; // beq 2 $zero _ElseBegin41_
	HD[1326] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[1327] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1328] = 32'b001011_00000000000000010101000011; // jump _IfExit41_
	HD[1329] = 32'b000101_00000_00010_0000000000000001; // li 2 1 / _ElseBegin41_
	HD[1330] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[1331] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[1332] = 32'b100111_10001_00000_00000_00001110000; // lcdwrite 17 112
	HD[1333] = 32'b100111_10010_00000_00000_00001110010; // lcdwrite 18 114
	HD[1334] = 32'b100111_10011_00000_00000_00001101111; // lcdwrite 19 111
	HD[1335] = 32'b100111_10100_00000_00000_00001100111; // lcdwrite 20 103
	HD[1336] = 32'b100111_10101_00000_00000_00001110010; // lcdwrite 21 114
	HD[1337] = 32'b100111_10110_00000_00000_00001100001; // lcdwrite 22 97
	HD[1338] = 32'b100111_10111_00000_00000_00001101101; // lcdwrite 23 109
	HD[1339] = 32'b100111_11000_00000_00000_00001100001; // lcdwrite 24 97
	HD[1340] = 32'b100111_11001_00000_00000_00001110011; // lcdwrite 25 115
	HD[1341] = 32'b100111_11010_00000_00000_00000100000; // lcdwrite 26 32
	HD[1342] = 32'b100111_11011_00000_00000_00000111110; // lcdwrite 27 62
	HD[1343] = 32'b100111_11100_00000_00000_00000100000; // lcdwrite 28 32
	HD[1344] = 32'b100111_11101_00000_00000_00000110001; // lcdwrite 29 49
	HD[1345] = 32'b100111_11110_00000_00000_00000110000; // lcdwrite 30 48
	HD[1346] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[1347] = 32'b001011_00000000000000010101010110; // jump _IfExit40_ / _IfExit41_
	HD[1348] = 32'b000101_00000_00010_0000000000000001; // li 2 1 / _ElseBegin40_
	HD[1349] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[1350] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[1351] = 32'b100111_10001_00000_00000_00001110000; // lcdwrite 17 112
	HD[1352] = 32'b100111_10010_00000_00000_00001110010; // lcdwrite 18 114
	HD[1353] = 32'b100111_10011_00000_00000_00001101111; // lcdwrite 19 111
	HD[1354] = 32'b100111_10100_00000_00000_00001100111; // lcdwrite 20 103
	HD[1355] = 32'b100111_10101_00000_00000_00001110010; // lcdwrite 21 114
	HD[1356] = 32'b100111_10110_00000_00000_00001100001; // lcdwrite 22 97
	HD[1357] = 32'b100111_10111_00000_00000_00001101101; // lcdwrite 23 109
	HD[1358] = 32'b100111_11000_00000_00000_00001100001; // lcdwrite 24 97
	HD[1359] = 32'b100111_11001_00000_00000_00001110011; // lcdwrite 25 115
	HD[1360] = 32'b100111_11010_00000_00000_00000100000; // lcdwrite 26 32
	HD[1361] = 32'b100111_11011_00000_00000_00000111100; // lcdwrite 27 60
	HD[1362] = 32'b100111_11100_00000_00000_00000100000; // lcdwrite 28 32
	HD[1363] = 32'b100111_11101_00000_00000_00000110000; // lcdwrite 29 48
	HD[1364] = 32'b100111_11110_00000_00000_00000100000; // lcdwrite 30 32
	HD[1365] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[1366] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2 / _IfExit40_
	HD[1367] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[1368] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1369] = 32'b000111_00010_00000_0000000000001111; // beq 2 $zero _IfExit42_
	HD[1370] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1371] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1372] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1373] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1374] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1375] = 32'b000101_00000_00010_0000000000000010; // li 2 2
	HD[1376] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1377] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1378] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1379] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1380] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1381] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1382] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[1383] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[1384] = 32'b001011_00000000000000010011111110; // jump _WhileBegin12_ / _IfExit42_
	HD[1385] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileExit12_ _WhileBegin13_
	HD[1386] = 32'b000001_10101_00011_0000000000000001; // lw 3 $fp 1
	HD[1387] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[1388] = 32'b000111_00010_00000_0000000010001111; // beq 2 $zero _WhileExit13_
	HD[1389] = 32'b000101_00000_00010_0000000000000010; // li 2 2
	HD[1390] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1391] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1392] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1393] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1394] = 32'b100111_10000_00000_00000_00001110000; // lcdwrite 16 112
	HD[1395] = 32'b100111_10001_00000_00000_00001100001; // lcdwrite 17 97
	HD[1396] = 32'b100111_10010_00000_00000_00001110010; // lcdwrite 18 114
	HD[1397] = 32'b100111_10011_00000_00000_00001100001; // lcdwrite 19 97
	HD[1398] = 32'b100111_10100_00000_00000_00000100000; // lcdwrite 20 32
	HD[1399] = 32'b100111_10101_00000_00000_00001110011; // lcdwrite 21 115
	HD[1400] = 32'b100111_10110_00000_00000_00001100101; // lcdwrite 22 101
	HD[1401] = 32'b100111_10111_00000_00000_00001110010; // lcdwrite 23 114
	HD[1402] = 32'b100111_11000_00000_00000_00000100000; // lcdwrite 24 32
	HD[1403] = 32'b100111_11001_00000_00000_00001100001; // lcdwrite 25 97
	HD[1404] = 32'b100111_11010_00000_00000_00001101100; // lcdwrite 26 108
	HD[1405] = 32'b100111_11011_00000_00000_00001101111; // lcdwrite 27 111
	HD[1406] = 32'b100111_11100_00000_00000_00001100011; // lcdwrite 28 99
	HD[1407] = 32'b100111_11101_00000_00000_00001100001; // lcdwrite 29 97
	HD[1408] = 32'b100111_11110_00000_00000_00001100100; // lcdwrite 30 100
	HD[1409] = 32'b100111_11111_00000_00000_00001101111; // lcdwrite 31 111
	HD[1410] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[1411] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[1412] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3
	HD[1413] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1414] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1415] = 32'b101000_00000000000000001001100110; // jal posicao_programa
	HD[1416] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1417] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[1418] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[1419] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1420] = 32'b000111_00010_00000_0000000000010100; // beq 2 $zero _ElseBegin43_
	HD[1421] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1422] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[1423] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[1424] = 32'b100111_10001_00000_00000_00001110000; // lcdwrite 17 112
	HD[1425] = 32'b100111_10010_00000_00000_00001110010; // lcdwrite 18 114
	HD[1426] = 32'b100111_10011_00000_00000_00001101111; // lcdwrite 19 111
	HD[1427] = 32'b100111_10100_00000_00000_00001100111; // lcdwrite 20 103
	HD[1428] = 32'b100111_10101_00000_00000_00000101110; // lcdwrite 21 46
	HD[1429] = 32'b100111_10110_00000_00000_00000100000; // lcdwrite 22 32
	HD[1430] = 32'b100111_10111_00000_00000_00001101001; // lcdwrite 23 105
	HD[1431] = 32'b100111_11000_00000_00000_00001101110; // lcdwrite 24 110
	HD[1432] = 32'b100111_11001_00000_00000_00001110110; // lcdwrite 25 118
	HD[1433] = 32'b100111_11010_00000_00000_00001100001; // lcdwrite 26 97
	HD[1434] = 32'b100111_11011_00000_00000_00001101100; // lcdwrite 27 108
	HD[1435] = 32'b100111_11100_00000_00000_00001101001; // lcdwrite 28 105
	HD[1436] = 32'b100111_11101_00000_00000_00001100100; // lcdwrite 29 100
	HD[1437] = 32'b100111_11110_00000_00000_00001101111; // lcdwrite 30 111
	HD[1438] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[1439] = 32'b001011_00000000000000010111101000; // jump _IfExit43_
	HD[1440] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3 / _ElseBegin43_
	HD[1441] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1442] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1443] = 32'b101000_00000000000000000111101000; // jal fila_existe_processo
	HD[1444] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1445] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[1446] = 32'b000001_00000_00011_0000000000010110; // lw 3 $global 22
	HD[1447] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1448] = 32'b000111_00010_00000_0000000000101110; // beq 2 $zero _ElseBegin44_
	HD[1449] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3
	HD[1450] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1451] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1452] = 32'b101000_00000000000000001000011111; // jal insere_processo_fila_pronto
	HD[1453] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1454] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[1455] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[1456] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1457] = 32'b100110_00000000000000000000000000; // lcdclean
	HD[1458] = 32'b000101_00000_00010_0000000000000101; // li 2 5
	HD[1459] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1460] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1461] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1462] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1463] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3
	HD[1464] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1465] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[1466] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1467] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[1468] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1469] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1470] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[1471] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1472] = 32'b100111_10000_00000_00000_00001101001; // lcdwrite 16 105
	HD[1473] = 32'b100111_10001_00000_00000_00001101110; // lcdwrite 17 110
	HD[1474] = 32'b100111_10010_00000_00000_00001110011; // lcdwrite 18 115
	HD[1475] = 32'b100111_10011_00000_00000_00001100101; // lcdwrite 19 101
	HD[1476] = 32'b100111_10100_00000_00000_00001110010; // lcdwrite 20 114
	HD[1477] = 32'b100111_10101_00000_00000_00001101001; // lcdwrite 21 105
	HD[1478] = 32'b100111_10110_00000_00000_00001100100; // lcdwrite 22 100
	HD[1479] = 32'b100111_10111_00000_00000_00001101111; // lcdwrite 23 111
	HD[1480] = 32'b100111_11001_00000_00000_00001101110; // lcdwrite 25 110
	HD[1481] = 32'b100111_11010_00000_00000_00001100001; // lcdwrite 26 97
	HD[1482] = 32'b100111_11100_00000_00000_00001100110; // lcdwrite 28 102
	HD[1483] = 32'b100111_11101_00000_00000_00001101001; // lcdwrite 29 105
	HD[1484] = 32'b100111_11110_00000_00000_00001101100; // lcdwrite 30 108
	HD[1485] = 32'b100111_11111_00000_00000_00001100001; // lcdwrite 31 97
	HD[1486] = 32'b000101_00000_00010_0000000000000010; // li 2 2
	HD[1487] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1488] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1489] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1490] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1491] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1492] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1493] = 32'b001011_00000000000000010111101000; // jump _IfExit44_
	HD[1494] = 32'b000101_00000_00010_0000000000000001; // li 2 1 / _ElseBegin44_
	HD[1495] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[1496] = 32'b100111_10000_00000_00000_00001110000; // lcdwrite 16 112
	HD[1497] = 32'b100111_10001_00000_00000_00001110010; // lcdwrite 17 114
	HD[1498] = 32'b100111_10010_00000_00000_00001101111; // lcdwrite 18 111
	HD[1499] = 32'b100111_10011_00000_00000_00001100011; // lcdwrite 19 99
	HD[1500] = 32'b100111_10100_00000_00000_00000101110; // lcdwrite 20 46
	HD[1501] = 32'b100111_10101_00000_00000_00000100000; // lcdwrite 21 32
	HD[1502] = 32'b100111_10110_00000_00000_00001101010; // lcdwrite 22 106
	HD[1503] = 32'b100111_10111_00000_00000_00001100001; // lcdwrite 23 97
	HD[1504] = 32'b100111_11000_00000_00000_00000100000; // lcdwrite 24 32
	HD[1505] = 32'b100111_11001_00000_00000_00001100001; // lcdwrite 25 97
	HD[1506] = 32'b100111_11010_00000_00000_00001101100; // lcdwrite 26 108
	HD[1507] = 32'b100111_11011_00000_00000_00001101111; // lcdwrite 27 111
	HD[1508] = 32'b100111_11100_00000_00000_00001100011; // lcdwrite 28 99
	HD[1509] = 32'b100111_11101_00000_00000_00001100001; // lcdwrite 29 97
	HD[1510] = 32'b100111_11110_00000_00000_00001100100; // lcdwrite 30 100
	HD[1511] = 32'b100111_11111_00000_00000_00001101111; // lcdwrite 31 111
	HD[1512] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2 / _IfExit44_ _IfExit43_
	HD[1513] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[1514] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1515] = 32'b000111_00010_00000_0000000000001111; // beq 2 $zero _IfExit45_
	HD[1516] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1517] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1518] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1519] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1520] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1521] = 32'b000101_00000_00010_0000000000000010; // li 2 2
	HD[1522] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1523] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1524] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1525] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1526] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1527] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1528] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[1529] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[1530] = 32'b001011_00000000000000010101101001; // jump _WhileBegin13_ / _IfExit45_
	HD[1531] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _WhileExit13_ _IfExit39_
	HD[1532] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[1533] = 32'b001111_10110_10111_0000000000000000; // push $ra / menu_opt0_executar_prog
	HD[1534] = 32'b100111_00000_00000_00000_00000100000; // lcdwrite 0 32
	HD[1535] = 32'b100111_00001_00000_00000_00000100000; // lcdwrite 1 32
	HD[1536] = 32'b100111_00010_00000_00000_00001000001; // lcdwrite 2 65
	HD[1537] = 32'b100111_00011_00000_00000_00001110100; // lcdwrite 3 116
	HD[1538] = 32'b100111_00100_00000_00000_00001101001; // lcdwrite 4 105
	HD[1539] = 32'b100111_00101_00000_00000_00001110110; // lcdwrite 5 118
	HD[1540] = 32'b100111_00110_00000_00000_00001100001; // lcdwrite 6 97
	HD[1541] = 32'b100111_00111_00000_00000_00001110010; // lcdwrite 7 114
	HD[1542] = 32'b100111_01000_00000_00000_00000100000; // lcdwrite 8 32
	HD[1543] = 32'b100111_01001_00000_00000_00000100000; // lcdwrite 9 32
	HD[1544] = 32'b100111_01010_00000_00000_00001101101; // lcdwrite 10 109
	HD[1545] = 32'b100111_01011_00000_00000_00001101111; // lcdwrite 11 111
	HD[1546] = 32'b100111_01100_00000_00000_00001100100; // lcdwrite 12 100
	HD[1547] = 32'b100111_01101_00000_00000_00001101111; // lcdwrite 13 111
	HD[1548] = 32'b100111_01110_00000_00000_00000100000; // lcdwrite 14 32
	HD[1549] = 32'b100111_01111_00000_00000_00000100000; // lcdwrite 15 32
	HD[1550] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[1551] = 32'b100111_10001_00000_00000_00001110000; // lcdwrite 17 112
	HD[1552] = 32'b100111_10010_00000_00000_00001110010; // lcdwrite 18 114
	HD[1553] = 32'b100111_10011_00000_00000_00001100101; // lcdwrite 19 101
	HD[1554] = 32'b100111_10100_00000_00000_00001100101; // lcdwrite 20 101
	HD[1555] = 32'b100111_10101_00000_00000_00001101101; // lcdwrite 21 109
	HD[1556] = 32'b100111_10110_00000_00000_00001110000; // lcdwrite 22 112
	HD[1557] = 32'b100111_10111_00000_00000_00001110100; // lcdwrite 23 116
	HD[1558] = 32'b100111_11000_00000_00000_00001101001; // lcdwrite 24 105
	HD[1559] = 32'b100111_11001_00000_00000_00001110110; // lcdwrite 25 118
	HD[1560] = 32'b100111_11010_00000_00000_00001101111; // lcdwrite 26 111
	HD[1561] = 32'b100111_11011_00000_00000_00000111111; // lcdwrite 27 63
	HD[1562] = 32'b100111_11100_00000_00000_00000100000; // lcdwrite 28 32
	HD[1563] = 32'b100111_11101_00000_00000_00001111001; // lcdwrite 29 121
	HD[1564] = 32'b100111_11110_00000_00000_00000111110; // lcdwrite 30 62
	HD[1565] = 32'b100111_11111_00000_00000_00000110000; // lcdwrite 31 48
	HD[1566] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[1567] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[1568] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _WhileBegin14_
	HD[1569] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1570] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[1571] = 32'b000111_00010_00000_0000000000000100; // beq 2 $zero _WhileExit14_
	HD[1572] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[1573] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[1574] = 32'b001011_00000000000000011000100000; // jump _WhileBegin14_
	HD[1575] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2 / _WhileExit14_
	HD[1576] = 32'b101000_00000000000000010011110101; // jal seleciona_programas
	HD[1577] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[1578] = 32'b100110_00000000000000000000000000; // lcdclean
	HD[1579] = 32'b100111_00001_00000_00000_00001001001; // lcdwrite 1 73
	HD[1580] = 32'b100111_00010_00000_00000_00001101110; // lcdwrite 2 110
	HD[1581] = 32'b100111_00011_00000_00000_00001101001; // lcdwrite 3 105
	HD[1582] = 32'b100111_00100_00000_00000_00001100011; // lcdwrite 4 99
	HD[1583] = 32'b100111_00101_00000_00000_00001101001; // lcdwrite 5 105
	HD[1584] = 32'b100111_00110_00000_00000_00001100001; // lcdwrite 6 97
	HD[1585] = 32'b100111_00111_00000_00000_00001101110; // lcdwrite 7 110
	HD[1586] = 32'b100111_01000_00000_00000_00001100100; // lcdwrite 8 100
	HD[1587] = 32'b100111_01001_00000_00000_00001101111; // lcdwrite 9 111
	HD[1588] = 32'b100111_01011_00000_00000_00001100101; // lcdwrite 11 101
	HD[1589] = 32'b100111_01100_00000_00000_00001111000; // lcdwrite 12 120
	HD[1590] = 32'b100111_01101_00000_00000_00001100101; // lcdwrite 13 101
	HD[1591] = 32'b100111_01110_00000_00000_00001100011; // lcdwrite 14 99
	HD[1592] = 32'b100111_10001_00000_00000_00000111110; // lcdwrite 17 62
	HD[1593] = 32'b100111_10010_00000_00000_00000111110; // lcdwrite 18 62
	HD[1594] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1595] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1596] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[1597] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1598] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1599] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1600] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[1601] = 32'b100111_10111_00000_00000_00000111110; // lcdwrite 23 62
	HD[1602] = 32'b100111_11000_00000_00000_00000111110; // lcdwrite 24 62
	HD[1603] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1604] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1605] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[1606] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1607] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1608] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1609] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[1610] = 32'b100111_11101_00000_00000_00000111110; // lcdwrite 29 62
	HD[1611] = 32'b100111_11110_00000_00000_00000111110; // lcdwrite 30 62
	HD[1612] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1613] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1614] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[1615] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1616] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1617] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1618] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[1619] = 32'b000001_00000_00010_0000000000001000; // lw 2 $global 8
	HD[1620] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[1621] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1622] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin46_
	HD[1623] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[1624] = 32'b101000_00000000000000001110110111; // jal executa_processos
	HD[1625] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[1626] = 32'b001011_00000000000000011001100110; // jump _IfExit46_
	HD[1627] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _ElseBegin46_
	HD[1628] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1629] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1630] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin47_
	HD[1631] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[1632] = 32'b101000_00000000000000001110110111; // jal executa_processos
	HD[1633] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[1634] = 32'b001011_00000000000000011001100110; // jump _IfExit47_
	HD[1635] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2 / _ElseBegin47_
	HD[1636] = 32'b101000_00000000000000010000000101; // jal executa_processos_preemptivo
	HD[1637] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[1638] = 32'b100111_00000_00000_00000_00000100000; // lcdwrite 0 32 / _IfExit47_ _IfExit46_
	HD[1639] = 32'b100111_00001_00000_00000_00000101101; // lcdwrite 1 45
	HD[1640] = 32'b100111_00010_00000_00000_00000101101; // lcdwrite 2 45
	HD[1641] = 32'b100111_00011_00000_00000_00001010000; // lcdwrite 3 80
	HD[1642] = 32'b100111_00100_00000_00000_00001110010; // lcdwrite 4 114
	HD[1643] = 32'b100111_00101_00000_00000_00001101111; // lcdwrite 5 111
	HD[1644] = 32'b100111_00110_00000_00000_00001100011; // lcdwrite 6 99
	HD[1645] = 32'b100111_00111_00000_00000_00001100101; // lcdwrite 7 101
	HD[1646] = 32'b100111_01000_00000_00000_00001110011; // lcdwrite 8 115
	HD[1647] = 32'b100111_01001_00000_00000_00001110011; // lcdwrite 9 115
	HD[1648] = 32'b100111_01010_00000_00000_00001101111; // lcdwrite 10 111
	HD[1649] = 32'b100111_01011_00000_00000_00001110011; // lcdwrite 11 115
	HD[1650] = 32'b100111_01100_00000_00000_00000101101; // lcdwrite 12 45
	HD[1651] = 32'b100111_01101_00000_00000_00000101101; // lcdwrite 13 45
	HD[1652] = 32'b100111_01110_00000_00000_00000101101; // lcdwrite 14 45
	HD[1653] = 32'b100111_01111_00000_00000_00000100000; // lcdwrite 15 32
	HD[1654] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[1655] = 32'b100111_10001_00000_00000_00000101101; // lcdwrite 17 45
	HD[1656] = 32'b100111_10010_00000_00000_00000101101; // lcdwrite 18 45
	HD[1657] = 32'b100111_10011_00000_00000_00001000110; // lcdwrite 19 70
	HD[1658] = 32'b100111_10100_00000_00000_00001101001; // lcdwrite 20 105
	HD[1659] = 32'b100111_10101_00000_00000_00001101110; // lcdwrite 21 110
	HD[1660] = 32'b100111_10110_00000_00000_00001100001; // lcdwrite 22 97
	HD[1661] = 32'b100111_10111_00000_00000_00001101100; // lcdwrite 23 108
	HD[1662] = 32'b100111_11000_00000_00000_00001101001; // lcdwrite 24 105
	HD[1663] = 32'b100111_11001_00000_00000_00001111010; // lcdwrite 25 122
	HD[1664] = 32'b100111_11010_00000_00000_00001100001; // lcdwrite 26 97
	HD[1665] = 32'b100111_11011_00000_00000_00001100100; // lcdwrite 27 100
	HD[1666] = 32'b100111_11100_00000_00000_00001101111; // lcdwrite 28 111
	HD[1667] = 32'b100111_11101_00000_00000_00001110011; // lcdwrite 29 115
	HD[1668] = 32'b100111_11110_00000_00000_00000101101; // lcdwrite 30 45
	HD[1669] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[1670] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[1671] = 32'b001010_00010_00000_0000000000000000; // out 2
	HD[1672] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[1673] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[1674] = 32'b001111_10110_10111_0000000000000000; // push $ra / menu_opt1_escrever_prog
	HD[1675] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[1676] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[1677] = 32'b100111_00000_00000_00000_00001000100; // lcdwrite 0 68
	HD[1678] = 32'b100111_00001_00000_00000_00001100101; // lcdwrite 1 101
	HD[1679] = 32'b100111_00010_00000_00000_00001110100; // lcdwrite 2 116
	HD[1680] = 32'b100111_00011_00000_00000_00001100101; // lcdwrite 3 101
	HD[1681] = 32'b100111_00100_00000_00000_00001110010; // lcdwrite 4 114
	HD[1682] = 32'b100111_00101_00000_00000_00001101101; // lcdwrite 5 109
	HD[1683] = 32'b100111_00110_00000_00000_00001101001; // lcdwrite 6 105
	HD[1684] = 32'b100111_00111_00000_00000_00001101110; // lcdwrite 7 110
	HD[1685] = 32'b100111_01000_00000_00000_00001100101; // lcdwrite 8 101
	HD[1686] = 32'b100111_01001_00000_00000_00000100000; // lcdwrite 9 32
	HD[1687] = 32'b100111_01010_00000_00000_00001110101; // lcdwrite 10 117
	HD[1688] = 32'b100111_01011_00000_00000_00001101101; // lcdwrite 11 109
	HD[1689] = 32'b100111_01100_00000_00000_00000100000; // lcdwrite 12 32
	HD[1690] = 32'b100111_01101_00000_00000_00001001001; // lcdwrite 13 73
	HD[1691] = 32'b100111_01110_00000_00000_00001000100; // lcdwrite 14 68
	HD[1692] = 32'b100111_01111_00000_00000_00000100000; // lcdwrite 15 32
	HD[1693] = 32'b100111_10000_00000_00000_00001110000; // lcdwrite 16 112
	HD[1694] = 32'b100111_10001_00000_00000_00001100001; // lcdwrite 17 97
	HD[1695] = 32'b100111_10010_00000_00000_00001110010; // lcdwrite 18 114
	HD[1696] = 32'b100111_10011_00000_00000_00001100001; // lcdwrite 19 97
	HD[1697] = 32'b100111_10100_00000_00000_00000100000; // lcdwrite 20 32
	HD[1698] = 32'b100111_10101_00000_00000_00001101111; // lcdwrite 21 111
	HD[1699] = 32'b100111_10110_00000_00000_00000100000; // lcdwrite 22 32
	HD[1700] = 32'b100111_10111_00000_00000_00001110000; // lcdwrite 23 112
	HD[1701] = 32'b100111_11000_00000_00000_00001110010; // lcdwrite 24 114
	HD[1702] = 32'b100111_11001_00000_00000_00001101111; // lcdwrite 25 111
	HD[1703] = 32'b100111_11010_00000_00000_00001100111; // lcdwrite 26 103
	HD[1704] = 32'b100111_11011_00000_00000_00001110010; // lcdwrite 27 114
	HD[1705] = 32'b100111_11100_00000_00000_00001100001; // lcdwrite 28 97
	HD[1706] = 32'b100111_11101_00000_00000_00001101101; // lcdwrite 29 109
	HD[1707] = 32'b100111_11110_00000_00000_00001100001; // lcdwrite 30 97
	HD[1708] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[1709] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[1710] = 32'b000101_00000_00011_0000001111101000; // li 3 1000
	HD[1711] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1712] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1713] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1714] = 32'b101000_00000000000000000001011010; // jal mod
	HD[1715] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1716] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[1717] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[1718] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[1719] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1720] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
	HD[1721] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[1722] = 32'b000111_00010_00000_0000000000001001; // beq 2 $zero _ElseBegin48_
	HD[1723] = 32'b000101_00000_00010_0000000000000110; // li 2 6
	HD[1724] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1725] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1726] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1727] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1728] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1729] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[1730] = 32'b001011_00000000000000011101010011; // jump _IfExit48_
	HD[1731] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _ElseBegin48_
	HD[1732] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1733] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1734] = 32'b101000_00000000000000001001100110; // jal posicao_programa
	HD[1735] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1736] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[1737] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[1738] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1739] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[1740] = 32'b000111_00010_00000_0000000000010101; // beq 2 $zero _ElseBegin49_
	HD[1741] = 32'b000101_00000_00010_0000000000000101; // li 2 5
	HD[1742] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1743] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1744] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1745] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1746] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[1747] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1748] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[1749] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1750] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[1751] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1752] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1753] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[1754] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1755] = 32'b000101_00000_00010_0000000000000111; // li 2 7
	HD[1756] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1757] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1758] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1759] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1760] = 32'b001011_00000000000000011101010011; // jump _IfExit49_
	HD[1761] = 32'b100110_00000000000000000000000000; // lcdclean / _ElseBegin49_
	HD[1762] = 32'b100111_00000_00000_00000_00001000100; // lcdwrite 0 68
	HD[1763] = 32'b100111_00001_00000_00000_00001100101; // lcdwrite 1 101
	HD[1764] = 32'b100111_00010_00000_00000_00001110100; // lcdwrite 2 116
	HD[1765] = 32'b100111_00011_00000_00000_00001100101; // lcdwrite 3 101
	HD[1766] = 32'b100111_00100_00000_00000_00001110010; // lcdwrite 4 114
	HD[1767] = 32'b100111_00101_00000_00000_00001101101; // lcdwrite 5 109
	HD[1768] = 32'b100111_00110_00000_00000_00001101001; // lcdwrite 6 105
	HD[1769] = 32'b100111_00111_00000_00000_00001101110; // lcdwrite 7 110
	HD[1770] = 32'b100111_01000_00000_00000_00001100101; // lcdwrite 8 101
	HD[1771] = 32'b100111_01010_00000_00000_00001101111; // lcdwrite 10 111
	HD[1772] = 32'b100111_01100_00000_00000_00001010100; // lcdwrite 12 84
	HD[1773] = 32'b100111_01101_00000_00000_00001100001; // lcdwrite 13 97
	HD[1774] = 32'b100111_01110_00000_00000_00001101101; // lcdwrite 14 109
	HD[1775] = 32'b100111_10010_00000_00000_00001100100; // lcdwrite 18 100
	HD[1776] = 32'b100111_10011_00000_00000_00001101111; // lcdwrite 19 111
	HD[1777] = 32'b100111_10101_00000_00000_00001110000; // lcdwrite 21 112
	HD[1778] = 32'b100111_10110_00000_00000_00001110010; // lcdwrite 22 114
	HD[1779] = 32'b100111_10111_00000_00000_00001101111; // lcdwrite 23 111
	HD[1780] = 32'b100111_11000_00000_00000_00001100111; // lcdwrite 24 103
	HD[1781] = 32'b100111_11001_00000_00000_00001110010; // lcdwrite 25 114
	HD[1782] = 32'b100111_11010_00000_00000_00001100001; // lcdwrite 26 97
	HD[1783] = 32'b100111_11011_00000_00000_00001101101; // lcdwrite 27 109
	HD[1784] = 32'b100111_11100_00000_00000_00001100001; // lcdwrite 28 97
	HD[1785] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[1786] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[1787] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[1788] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1789] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
	HD[1790] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[1791] = 32'b000111_00010_00000_0000000000010100; // beq 2 $zero _ElseBegin50_
	HD[1792] = 32'b100111_10000_00000_00000_00001010100; // lcdwrite 16 84
	HD[1793] = 32'b100111_10001_00000_00000_00001100001; // lcdwrite 17 97
	HD[1794] = 32'b100111_10010_00000_00000_00001101101; // lcdwrite 18 109
	HD[1795] = 32'b100111_10011_00000_00000_00000100000; // lcdwrite 19 32
	HD[1796] = 32'b100111_10100_00000_00000_00001100100; // lcdwrite 20 100
	HD[1797] = 32'b100111_10101_00000_00000_00001100101; // lcdwrite 21 101
	HD[1798] = 32'b100111_10110_00000_00000_00001110110; // lcdwrite 22 118
	HD[1799] = 32'b100111_10111_00000_00000_00001100101; // lcdwrite 23 101
	HD[1800] = 32'b100111_11000_00000_00000_00000100000; // lcdwrite 24 32
	HD[1801] = 32'b100111_11001_00000_00000_00001110011; // lcdwrite 25 115
	HD[1802] = 32'b100111_11010_00000_00000_00001100101; // lcdwrite 26 101
	HD[1803] = 32'b100111_11011_00000_00000_00001110010; // lcdwrite 27 114
	HD[1804] = 32'b100111_11100_00000_00000_00000100000; // lcdwrite 28 32
	HD[1805] = 32'b100111_11101_00000_00000_00000111110; // lcdwrite 29 62
	HD[1806] = 32'b100111_11110_00000_00000_00000100000; // lcdwrite 30 32
	HD[1807] = 32'b100111_11111_00000_00000_00000110000; // lcdwrite 31 48
	HD[1808] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1809] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[1810] = 32'b001011_00000000000000011101010011; // jump _IfExit50_
	HD[1811] = 32'b100110_00000000000000000000000000; // lcdclean / _ElseBegin50_
	HD[1812] = 32'b100111_00000_00000_00000_00001001001; // lcdwrite 0 73
	HD[1813] = 32'b100111_00001_00000_00000_00001101110; // lcdwrite 1 110
	HD[1814] = 32'b100111_00010_00000_00000_00001110011; // lcdwrite 2 115
	HD[1815] = 32'b100111_00011_00000_00000_00001101001; // lcdwrite 3 105
	HD[1816] = 32'b100111_00100_00000_00000_00001110010; // lcdwrite 4 114
	HD[1817] = 32'b100111_00101_00000_00000_00001100001; // lcdwrite 5 97
	HD[1818] = 32'b100111_00110_00000_00000_00000111010; // lcdwrite 6 58
	HD[1819] = 32'b100111_01000_00000_00000_00001101001; // lcdwrite 8 105
	HD[1820] = 32'b100111_01001_00000_00000_00001101110; // lcdwrite 9 110
	HD[1821] = 32'b100111_01010_00000_00000_00001110011; // lcdwrite 10 115
	HD[1822] = 32'b100111_01011_00000_00000_00001110100; // lcdwrite 11 116
	HD[1823] = 32'b100111_10000_00000_00000_00001100100; // lcdwrite 16 100
	HD[1824] = 32'b100111_10001_00000_00000_00001101111; // lcdwrite 17 111
	HD[1825] = 32'b100111_10011_00000_00000_00001010000; // lcdwrite 19 80
	HD[1826] = 32'b100111_10100_00000_00000_00001110010; // lcdwrite 20 114
	HD[1827] = 32'b100111_10101_00000_00000_00001101111; // lcdwrite 21 111
	HD[1828] = 32'b100111_10110_00000_00000_00001100111; // lcdwrite 22 103
	HD[1829] = 32'b100111_10111_00000_00000_00001110010; // lcdwrite 23 114
	HD[1830] = 32'b100111_11000_00000_00000_00001100001; // lcdwrite 24 97
	HD[1831] = 32'b100111_11001_00000_00000_00001101101; // lcdwrite 25 109
	HD[1832] = 32'b100111_11010_00000_00000_00001100001; // lcdwrite 26 97
	HD[1833] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[1834] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[1835] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[1836] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1837] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[1838] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1839] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1840] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[1841] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1842] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[1843] = 32'b000001_10101_00011_0000000000000010; // lw 3 $fp 2
	HD[1844] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1845] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1846] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1847] = 32'b101000_00000000000000001011111111; // jal cria_programa
	HD[1848] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1849] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[1850] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1851] = 32'b100110_00000000000000000000000000; // lcdclean
	HD[1852] = 32'b000101_00000_00010_0000000000000101; // li 2 5
	HD[1853] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1854] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1855] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1856] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1857] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[1858] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1859] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[1860] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1861] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[1862] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1863] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1864] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[1865] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1866] = 32'b100111_10011_00000_00000_00001100110; // lcdwrite 19 102
	HD[1867] = 32'b100111_10100_00000_00000_00001101111; // lcdwrite 20 111
	HD[1868] = 32'b100111_10101_00000_00000_00001101001; // lcdwrite 21 105
	HD[1869] = 32'b100111_10111_00000_00000_00001100011; // lcdwrite 23 99
	HD[1870] = 32'b100111_11000_00000_00000_00001110010; // lcdwrite 24 114
	HD[1871] = 32'b100111_11001_00000_00000_00001101001; // lcdwrite 25 105
	HD[1872] = 32'b100111_11010_00000_00000_00001100001; // lcdwrite 26 97
	HD[1873] = 32'b100111_11011_00000_00000_00001100100; // lcdwrite 27 100
	HD[1874] = 32'b100111_11100_00000_00000_00001101111; // lcdwrite 28 111
	HD[1875] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3 / _IfExit50_ _IfExit49_ _IfExit48_
	HD[1876] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[1877] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1878] = 32'b000111_00010_00000_0000000000001111; // beq 2 $zero _IfExit51_
	HD[1879] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1880] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1881] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1882] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1883] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1884] = 32'b000101_00000_00010_0000000000000100; // li 2 4
	HD[1885] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1886] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1887] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1888] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1889] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[1890] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1891] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[1892] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[1893] = 32'b000101_00000_00010_0000000000000000; // li 2 0 / _IfExit51_
	HD[1894] = 32'b001010_00010_00000_0000000000000000; // out 2
	HD[1895] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[1896] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[1897] = 32'b001111_10110_10111_0000000000000000; // push $ra / menu_opt2_renomear_prog
	HD[1898] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[1899] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[1900] = 32'b000101_00000_00010_0000000000000010; // li 2 2
	HD[1901] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1902] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1903] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1904] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1905] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[1906] = 32'b100111_10001_00000_00000_00001100001; // lcdwrite 17 97
	HD[1907] = 32'b100111_10010_00000_00000_00000100000; // lcdwrite 18 32
	HD[1908] = 32'b100111_10011_00000_00000_00001110011; // lcdwrite 19 115
	HD[1909] = 32'b100111_10100_00000_00000_00001100101; // lcdwrite 20 101
	HD[1910] = 32'b100111_10101_00000_00000_00001110010; // lcdwrite 21 114
	HD[1911] = 32'b100111_10110_00000_00000_00000100000; // lcdwrite 22 32
	HD[1912] = 32'b100111_10111_00000_00000_00001110010; // lcdwrite 23 114
	HD[1913] = 32'b100111_11000_00000_00000_00001100101; // lcdwrite 24 101
	HD[1914] = 32'b100111_11001_00000_00000_00001101110; // lcdwrite 25 110
	HD[1915] = 32'b100111_11010_00000_00000_00001101111; // lcdwrite 26 111
	HD[1916] = 32'b100111_11011_00000_00000_00001101101; // lcdwrite 27 109
	HD[1917] = 32'b100111_11100_00000_00000_00001100101; // lcdwrite 28 101
	HD[1918] = 32'b100111_11101_00000_00000_00001100001; // lcdwrite 29 97
	HD[1919] = 32'b100111_11110_00000_00000_00001100100; // lcdwrite 30 100
	HD[1920] = 32'b100111_11111_00000_00000_00001101111; // lcdwrite 31 111
	HD[1921] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[1922] = 32'b000101_00000_00011_0000001111101000; // li 3 1000
	HD[1923] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1924] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1925] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1926] = 32'b101000_00000000000000000001011010; // jal mod
	HD[1927] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1928] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[1929] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[1930] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[1931] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1932] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
	HD[1933] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[1934] = 32'b000111_00010_00000_0000000000000100; // beq 2 $zero _ElseBegin52_
	HD[1935] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[1936] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[1937] = 32'b001011_00000000000000100000101011; // jump _IfExit52_
	HD[1938] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _ElseBegin52_
	HD[1939] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1940] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1941] = 32'b101000_00000000000000001001100110; // jal posicao_programa
	HD[1942] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1943] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[1944] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[1945] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[1946] = 32'b000111_00010_00000_0000000000010101; // beq 2 $zero _ElseBegin53_
	HD[1947] = 32'b000101_00000_00010_0000000000000011; // li 2 3
	HD[1948] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1949] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1950] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1951] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1952] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[1953] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[1954] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[1955] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1956] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[1957] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[1958] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1959] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[1960] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1961] = 32'b000101_00000_00010_0000000000000100; // li 2 4
	HD[1962] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[1963] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[1964] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[1965] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[1966] = 32'b001011_00000000000000100000101011; // jump _IfExit53_
	HD[1967] = 32'b100111_00000_00000_00000_00000100000; // lcdwrite 0 32 / _ElseBegin53_
	HD[1968] = 32'b100111_00001_00000_00000_00001000100; // lcdwrite 1 68
	HD[1969] = 32'b100111_00010_00000_00000_00001100101; // lcdwrite 2 101
	HD[1970] = 32'b100111_00011_00000_00000_00001100110; // lcdwrite 3 102
	HD[1971] = 32'b100111_00100_00000_00000_00001101001; // lcdwrite 4 105
	HD[1972] = 32'b100111_00101_00000_00000_00001101110; // lcdwrite 5 110
	HD[1973] = 32'b100111_00110_00000_00000_00001100001; // lcdwrite 6 97
	HD[1974] = 32'b100111_00111_00000_00000_00000100000; // lcdwrite 7 32
	HD[1975] = 32'b100111_01000_00000_00000_00001110101; // lcdwrite 8 117
	HD[1976] = 32'b100111_01001_00000_00000_00001101101; // lcdwrite 9 109
	HD[1977] = 32'b100111_01010_00000_00000_00000100000; // lcdwrite 10 32
	HD[1978] = 32'b100111_01011_00000_00000_00001101110; // lcdwrite 11 110
	HD[1979] = 32'b100111_01100_00000_00000_00001101111; // lcdwrite 12 111
	HD[1980] = 32'b100111_01101_00000_00000_00001110110; // lcdwrite 13 118
	HD[1981] = 32'b100111_01110_00000_00000_00001101111; // lcdwrite 14 111
	HD[1982] = 32'b100111_01111_00000_00000_00000100000; // lcdwrite 15 32
	HD[1983] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[1984] = 32'b100111_10001_00000_00000_00001001001; // lcdwrite 17 73
	HD[1985] = 32'b100111_10010_00000_00000_00001100100; // lcdwrite 18 100
	HD[1986] = 32'b100111_10011_00000_00000_00001100101; // lcdwrite 19 101
	HD[1987] = 32'b100111_10100_00000_00000_00001101110; // lcdwrite 20 110
	HD[1988] = 32'b100111_10101_00000_00000_00001110100; // lcdwrite 21 116
	HD[1989] = 32'b100111_10110_00000_00000_00001101001; // lcdwrite 22 105
	HD[1990] = 32'b100111_10111_00000_00000_00001100110; // lcdwrite 23 102
	HD[1991] = 32'b100111_11000_00000_00000_00001101001; // lcdwrite 24 105
	HD[1992] = 32'b100111_11001_00000_00000_00001100011; // lcdwrite 25 99
	HD[1993] = 32'b100111_11010_00000_00000_00001100001; // lcdwrite 26 97
	HD[1994] = 32'b100111_11011_00000_00000_00001100100; // lcdwrite 27 100
	HD[1995] = 32'b100111_11100_00000_00000_00001101111; // lcdwrite 28 111
	HD[1996] = 32'b100111_11101_00000_00000_00001110010; // lcdwrite 29 114
	HD[1997] = 32'b100111_11110_00000_00000_00000100000; // lcdwrite 30 32
	HD[1998] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[1999] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[2000] = 32'b000101_00000_00011_0000001111101000; // li 3 1000
	HD[2001] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2002] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2003] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2004] = 32'b101000_00000000000000000001011010; // jal mod
	HD[2005] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2006] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[2007] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[2008] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[2009] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2010] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
	HD[2011] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[2012] = 32'b000111_00010_00000_0000000000000100; // beq 2 $zero _ElseBegin54_
	HD[2013] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2014] = 32'b000010_10101_00010_0000000000000011; // sw 2 $fp 3
	HD[2015] = 32'b001011_00000000000000100000101011; // jump _IfExit54_
	HD[2016] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2 / _ElseBegin54_
	HD[2017] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2018] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2019] = 32'b101000_00000000000000001001100110; // jal posicao_programa
	HD[2020] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2021] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[2022] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[2023] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2024] = 32'b000111_00010_00000_0000000000110000; // beq 2 $zero _ElseBegin55_
	HD[2025] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[2026] = 32'b000001_10101_00011_0000000000000010; // lw 3 $fp 2
	HD[2027] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2028] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2029] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2030] = 32'b101000_00000000000000001101100111; // jal renomear_programa
	HD[2031] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2032] = 32'b000101_00000_00010_0000000000000101; // li 2 5
	HD[2033] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2034] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2035] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2036] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2037] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[2038] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2039] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[2040] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2041] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[2042] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2043] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2044] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[2045] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2046] = 32'b100111_10000_00000_00000_00001110010; // lcdwrite 16 114
	HD[2047] = 32'b100111_10001_00000_00000_00001100101; // lcdwrite 17 101
	HD[2048] = 32'b100111_10010_00000_00000_00001101110; // lcdwrite 18 110
	HD[2049] = 32'b100111_10011_00000_00000_00001101111; // lcdwrite 19 111
	HD[2050] = 32'b100111_10100_00000_00000_00001101101; // lcdwrite 20 109
	HD[2051] = 32'b100111_10101_00000_00000_00001100101; // lcdwrite 21 101
	HD[2052] = 32'b100111_10110_00000_00000_00001100001; // lcdwrite 22 97
	HD[2053] = 32'b100111_10111_00000_00000_00001100100; // lcdwrite 23 100
	HD[2054] = 32'b100111_11000_00000_00000_00001101111; // lcdwrite 24 111
	HD[2055] = 32'b100111_11001_00000_00000_00000100000; // lcdwrite 25 32
	HD[2056] = 32'b100111_11010_00000_00000_00001110000; // lcdwrite 26 112
	HD[2057] = 32'b100111_11011_00000_00000_00000101111; // lcdwrite 27 47
	HD[2058] = 32'b100111_11100_00000_00000_00000100000; // lcdwrite 28 32
	HD[2059] = 32'b100111_11101_00000_00000_00000100000; // lcdwrite 29 32
	HD[2060] = 32'b100111_11110_00000_00000_00000100000; // lcdwrite 30 32
	HD[2061] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2062] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[2063] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[2064] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[2065] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2066] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[2067] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2068] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2069] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[2070] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2071] = 32'b001011_00000000000000100000101011; // jump _IfExit55_
	HD[2072] = 32'b000101_00000_00010_0000000000000101; // li 2 5 / _ElseBegin55_
	HD[2073] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2074] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2075] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2076] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2077] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[2078] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2079] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[2080] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2081] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[2082] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2083] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2084] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[2085] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2086] = 32'b000101_00000_00010_0000000000000111; // li 2 7
	HD[2087] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2088] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2089] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2090] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2091] = 32'b000001_10101_00010_0000000000000011; // lw 2 $fp 3 / _IfExit55_ _IfExit54_ _IfExit53_ _IfExit52_
	HD[2092] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[2093] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2094] = 32'b000111_00010_00000_0000000000010100; // beq 2 $zero _IfExit56_
	HD[2095] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2096] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2097] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2098] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2099] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2100] = 32'b000101_00000_00010_0000000000000110; // li 2 6
	HD[2101] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2102] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2103] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2104] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2105] = 32'b000101_00000_00010_0000000000000100; // li 2 4
	HD[2106] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2107] = 32'b000011_10101_10101_0000000000000100; // addi $fp $fp 4
	HD[2108] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2109] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2110] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2111] = 32'b000100_10101_10101_0000000000000100; // subi $fp $fp 4
	HD[2112] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2113] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2114] = 32'b000101_00000_00010_0000000000000000; // li 2 0 / _IfExit56_
	HD[2115] = 32'b001010_00010_00000_0000000000000000; // out 2
	HD[2116] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2117] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2118] = 32'b001111_10110_10111_0000000000000000; // push $ra / menu_opt3_deletar_prog
	HD[2119] = 32'b000101_00000_00010_0000000000000010; // li 2 2
	HD[2120] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2121] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2122] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2123] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2124] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2125] = 32'b100111_10001_00000_00000_00001100001; // lcdwrite 17 97
	HD[2126] = 32'b100111_10010_00000_00000_00000100000; // lcdwrite 18 32
	HD[2127] = 32'b100111_10011_00000_00000_00001110011; // lcdwrite 19 115
	HD[2128] = 32'b100111_10100_00000_00000_00001100101; // lcdwrite 20 101
	HD[2129] = 32'b100111_10101_00000_00000_00001110010; // lcdwrite 21 114
	HD[2130] = 32'b100111_10110_00000_00000_00000100000; // lcdwrite 22 32
	HD[2131] = 32'b100111_10111_00000_00000_00001100100; // lcdwrite 23 100
	HD[2132] = 32'b100111_11000_00000_00000_00001100101; // lcdwrite 24 101
	HD[2133] = 32'b100111_11001_00000_00000_00001101100; // lcdwrite 25 108
	HD[2134] = 32'b100111_11010_00000_00000_00001100101; // lcdwrite 26 101
	HD[2135] = 32'b100111_11011_00000_00000_00001110100; // lcdwrite 27 116
	HD[2136] = 32'b100111_11100_00000_00000_00001100001; // lcdwrite 28 97
	HD[2137] = 32'b100111_11101_00000_00000_00001100100; // lcdwrite 29 100
	HD[2138] = 32'b100111_11110_00000_00000_00001101111; // lcdwrite 30 111
	HD[2139] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2140] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[2141] = 32'b000101_00000_00011_0000001111101000; // li 3 1000
	HD[2142] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2143] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2144] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2145] = 32'b101000_00000000000000000001011010; // jal mod
	HD[2146] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2147] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[2148] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[2149] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[2150] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2151] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2152] = 32'b101000_00000000000000001101001101; // jal deleta_programa
	HD[2153] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2154] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[2155] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2156] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[2157] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2158] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
	HD[2159] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[2160] = 32'b000111_00010_00000_0000000000010101; // beq 2 $zero _ElseBegin57_
	HD[2161] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2162] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2163] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2164] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2165] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2166] = 32'b000101_00000_00010_0000000000000110; // li 2 6
	HD[2167] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2168] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2169] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2170] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2171] = 32'b000101_00000_00010_0000000000000100; // li 2 4
	HD[2172] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2173] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2174] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2175] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2176] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2177] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2178] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2179] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2180] = 32'b001011_00000000000000100010111011; // jump _IfExit57_
	HD[2181] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin57_
	HD[2182] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[2183] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2184] = 32'b000111_00010_00000_0000000000010101; // beq 2 $zero _ElseBegin58_
	HD[2185] = 32'b000101_00000_00010_0000000000000011; // li 2 3
	HD[2186] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2187] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2188] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2189] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2190] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[2191] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2192] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[2193] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2194] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[2195] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2196] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2197] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[2198] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2199] = 32'b000101_00000_00010_0000000000000100; // li 2 4
	HD[2200] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2201] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2202] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2203] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2204] = 32'b001011_00000000000000100010111011; // jump _IfExit58_
	HD[2205] = 32'b000101_00000_00010_0000000000000101; // li 2 5 / _ElseBegin58_
	HD[2206] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2207] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2208] = 32'b101000_00000000000000000010110011; // jal print_default_msg
	HD[2209] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2210] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[2211] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2212] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[2213] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2214] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[2215] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2216] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2217] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[2218] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2219] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2220] = 32'b100111_10001_00000_00000_00000100000; // lcdwrite 17 32
	HD[2221] = 32'b100111_10010_00000_00000_00001100110; // lcdwrite 18 102
	HD[2222] = 32'b100111_10011_00000_00000_00001101111; // lcdwrite 19 111
	HD[2223] = 32'b100111_10100_00000_00000_00001101001; // lcdwrite 20 105
	HD[2224] = 32'b100111_10101_00000_00000_00000100000; // lcdwrite 21 32
	HD[2225] = 32'b100111_10110_00000_00000_00001100100; // lcdwrite 22 100
	HD[2226] = 32'b100111_10111_00000_00000_00001100101; // lcdwrite 23 101
	HD[2227] = 32'b100111_11000_00000_00000_00001101100; // lcdwrite 24 108
	HD[2228] = 32'b100111_11001_00000_00000_00001100101; // lcdwrite 25 101
	HD[2229] = 32'b100111_11010_00000_00000_00001110100; // lcdwrite 26 116
	HD[2230] = 32'b100111_11011_00000_00000_00001100001; // lcdwrite 27 97
	HD[2231] = 32'b100111_11100_00000_00000_00001100100; // lcdwrite 28 100
	HD[2232] = 32'b100111_11101_00000_00000_00001101111; // lcdwrite 29 111
	HD[2233] = 32'b100111_11110_00000_00000_00000100000; // lcdwrite 30 32
	HD[2234] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2235] = 32'b000101_00000_00010_0000000000000000; // li 2 0 / _IfExit58_ _IfExit57_
	HD[2236] = 32'b001010_00010_00000_0000000000000000; // out 2
	HD[2237] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2238] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2239] = 32'b001111_10110_10111_0000000000000000; // push $ra / menu_opt4_listar_prog
	HD[2240] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2241] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2242] = 32'b000010_10101_00010_0000000000010001; // sw 2 $fp 17
	HD[2243] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin15_
	HD[2244] = 32'b000001_00000_00011_0000000000000000; // lw 3 $global 0
	HD[2245] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[2246] = 32'b000111_00010_00000_0000000000010111; // beq 2 $zero _WhileExit15_
	HD[2247] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[2248] = 32'b000011_10101_10101_0000000000010010; // addi $fp $fp 18
	HD[2249] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2250] = 32'b101000_00000000000000001110101001; // jal existe_programa_posicao
	HD[2251] = 32'b000100_10101_10101_0000000000010010; // subi $fp $fp 18
	HD[2252] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[2253] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[2254] = 32'b000000_00011_10101_00011_00000_000101; // add 3 3 $fp
	HD[2255] = 32'b000010_00011_00010_0000000000000001; // sw 2 3 1
	HD[2256] = 32'b000010_10101_00010_0000000000010000; // sw 2 $fp 16
	HD[2257] = 32'b000001_10101_00010_0000000000010000; // lw 2 $fp 16
	HD[2258] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[2259] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2260] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[2261] = 32'b000111_00010_00000_0000000000000100; // beq 2 $zero _IfExit59_
	HD[2262] = 32'b000001_10101_00010_0000000000010001; // lw 2 $fp 17
	HD[2263] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[2264] = 32'b000010_10101_00010_0000000000010001; // sw 2 $fp 17
	HD[2265] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _IfExit59_
	HD[2266] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[2267] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2268] = 32'b001011_00000000000000100011000011; // jump _WhileBegin15_
	HD[2269] = 32'b100110_00000000000000000000000000; // lcdclean / _WhileExit15_
	HD[2270] = 32'b100111_00001_00000_00000_00001010001; // lcdwrite 1 81
	HD[2271] = 32'b100111_00010_00000_00000_00001110100; // lcdwrite 2 116
	HD[2272] = 32'b100111_00011_00000_00000_00001100100; // lcdwrite 3 100
	HD[2273] = 32'b100111_00101_00000_00000_00001010000; // lcdwrite 5 80
	HD[2274] = 32'b100111_00110_00000_00000_00001110010; // lcdwrite 6 114
	HD[2275] = 32'b100111_00111_00000_00000_00001101111; // lcdwrite 7 111
	HD[2276] = 32'b100111_01000_00000_00000_00001100111; // lcdwrite 8 103
	HD[2277] = 32'b100111_01001_00000_00000_00001110011; // lcdwrite 9 115
	HD[2278] = 32'b100111_01010_00000_00000_00000111010; // lcdwrite 10 58
	HD[2279] = 32'b000001_10101_00010_0000000000010001; // lw 2 $fp 17
	HD[2280] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2281] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[2282] = 32'b000011_10101_10101_0000000000010010; // addi $fp $fp 18
	HD[2283] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[2284] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2285] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2286] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[2287] = 32'b000100_10101_10101_0000000000010010; // subi $fp $fp 18
	HD[2288] = 32'b100111_10011_00000_00000_00001101111; // lcdwrite 19 111
	HD[2289] = 32'b100111_10101_00000_00000_00001010000; // lcdwrite 21 80
	HD[2290] = 32'b100111_10110_00000_00000_00001110010; // lcdwrite 22 114
	HD[2291] = 32'b100111_10111_00000_00000_00001101111; // lcdwrite 23 111
	HD[2292] = 32'b100111_11000_00000_00000_00001100111; // lcdwrite 24 103
	HD[2293] = 32'b100111_11001_00000_00000_00000111010; // lcdwrite 25 58
	HD[2294] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2295] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2296] = 32'b000010_10101_00010_0000000000010001; // sw 2 $fp 17
	HD[2297] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin16_
	HD[2298] = 32'b000001_00000_00011_0000000000000000; // lw 3 $global 0
	HD[2299] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[2300] = 32'b000111_00010_00000_0000000000100101; // beq 2 $zero _WhileExit16_
	HD[2301] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[2302] = 32'b000000_00010_10101_00010_00000_000101; // add 2 2 $fp
	HD[2303] = 32'b000001_00010_00010_0000000000000001; // lw 2 2 1
	HD[2304] = 32'b000010_10101_00010_0000000000010000; // sw 2 $fp 16
	HD[2305] = 32'b000001_10101_00010_0000000000010000; // lw 2 $fp 16
	HD[2306] = 32'b000001_00000_00011_0000000000011001; // lw 3 $global 25
	HD[2307] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2308] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[2309] = 32'b000111_00010_00000_0000000000011000; // beq 2 $zero _IfExit60_
	HD[2310] = 32'b000001_10101_00010_0000000000010001; // lw 2 $fp 17
	HD[2311] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[2312] = 32'b000010_10101_00010_0000000000010001; // sw 2 $fp 17
	HD[2313] = 32'b000001_10101_00010_0000000000010001; // lw 2 $fp 17
	HD[2314] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[2315] = 32'b000101_00000_00100_0000000000000010; // li 4 2
	HD[2316] = 32'b000011_10101_10101_0000000000010010; // addi $fp $fp 18
	HD[2317] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[2318] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2319] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2320] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[2321] = 32'b000100_10101_10101_0000000000010010; // subi $fp $fp 18
	HD[2322] = 32'b000001_10101_00010_0000000000010000; // lw 2 $fp 16
	HD[2323] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[2324] = 32'b000101_00000_00100_0000000000001110; // li 4 14
	HD[2325] = 32'b000011_10101_10101_0000000000010010; // addi $fp $fp 18
	HD[2326] = 32'b000010_10101_00100_0000000000000010; // sw 4 $fp 2
	HD[2327] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2328] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2329] = 32'b101000_00000000000000000001100111; // jal print_value
	HD[2330] = 32'b000100_10101_10101_0000000000010010; // subi $fp $fp 18
	HD[2331] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2332] = 32'b001010_00010_00000_0000000000000000; // out 2
	HD[2333] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _IfExit60_
	HD[2334] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[2335] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2336] = 32'b001011_00000000000000100011111001; // jump _WhileBegin16_
	HD[2337] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _WhileExit16_
	HD[2338] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2339] = 32'b001111_10110_10111_0000000000000000; // push $ra / menu_opt5_reiniciar
	HD[2340] = 32'b100110_00000000000000000000000000; // lcdclean
	HD[2341] = 32'b100111_00010_00000_00000_00001010010; // lcdwrite 2 82
	HD[2342] = 32'b100111_00011_00000_00000_00001100101; // lcdwrite 3 101
	HD[2343] = 32'b100111_00100_00000_00000_00001101001; // lcdwrite 4 105
	HD[2344] = 32'b100111_00101_00000_00000_00001101110; // lcdwrite 5 110
	HD[2345] = 32'b100111_00110_00000_00000_00001101001; // lcdwrite 6 105
	HD[2346] = 32'b100111_00111_00000_00000_00001100011; // lcdwrite 7 99
	HD[2347] = 32'b100111_01000_00000_00000_00001101001; // lcdwrite 8 105
	HD[2348] = 32'b100111_01001_00000_00000_00001100001; // lcdwrite 9 97
	HD[2349] = 32'b100111_01010_00000_00000_00001101110; // lcdwrite 10 110
	HD[2350] = 32'b100111_01011_00000_00000_00001100100; // lcdwrite 11 100
	HD[2351] = 32'b100111_01100_00000_00000_00001101111; // lcdwrite 12 111
	HD[2352] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2353] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2354] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2355] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2356] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2357] = 32'b100111_10000_00000_00000_00000111110; // lcdwrite 16 62
	HD[2358] = 32'b100111_11111_00000_00000_00000111100; // lcdwrite 31 60
	HD[2359] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2360] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2361] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2362] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2363] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2364] = 32'b100111_10010_00000_00000_00000111110; // lcdwrite 18 62
	HD[2365] = 32'b100111_11101_00000_00000_00000111100; // lcdwrite 29 60
	HD[2366] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2367] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2368] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2369] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2370] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2371] = 32'b100111_10100_00000_00000_00000111110; // lcdwrite 20 62
	HD[2372] = 32'b100111_11011_00000_00000_00000111100; // lcdwrite 27 60
	HD[2373] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2374] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2375] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2376] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2377] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2378] = 32'b100111_10110_00000_00000_00000111110; // lcdwrite 22 62
	HD[2379] = 32'b100111_11001_00000_00000_00000111100; // lcdwrite 25 60
	HD[2380] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2381] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2382] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2383] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2384] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2385] = 32'b100110_00000000000000000000000000; // lcdclean
	HD[2386] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2387] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2388] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2389] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2390] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2391] = 32'b100001_00000000000000000000000000; // upbios
	HD[2392] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2393] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2394] = 32'b001111_10110_10111_0000000000000000; // push $ra / menu_opt6_desligar
	HD[2395] = 32'b100110_00000000000000000000000000; // lcdclean
	HD[2396] = 32'b100111_00011_00000_00000_00001000100; // lcdwrite 3 68
	HD[2397] = 32'b100111_00100_00000_00000_00001100101; // lcdwrite 4 101
	HD[2398] = 32'b100111_00101_00000_00000_00001110011; // lcdwrite 5 115
	HD[2399] = 32'b100111_00110_00000_00000_00001101100; // lcdwrite 6 108
	HD[2400] = 32'b100111_00111_00000_00000_00001101001; // lcdwrite 7 105
	HD[2401] = 32'b100111_01000_00000_00000_00001100111; // lcdwrite 8 103
	HD[2402] = 32'b100111_01001_00000_00000_00001100001; // lcdwrite 9 97
	HD[2403] = 32'b100111_01010_00000_00000_00001101110; // lcdwrite 10 110
	HD[2404] = 32'b100111_01011_00000_00000_00001100100; // lcdwrite 11 100
	HD[2405] = 32'b100111_01100_00000_00000_00001101111; // lcdwrite 12 111
	HD[2406] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2407] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2408] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2409] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2410] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2411] = 32'b100111_10000_00000_00000_00000111110; // lcdwrite 16 62
	HD[2412] = 32'b100111_11111_00000_00000_00000111100; // lcdwrite 31 60
	HD[2413] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2414] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2415] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2416] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2417] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2418] = 32'b100111_10010_00000_00000_00000111110; // lcdwrite 18 62
	HD[2419] = 32'b100111_11101_00000_00000_00000111100; // lcdwrite 29 60
	HD[2420] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2421] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2422] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2423] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2424] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2425] = 32'b100111_10100_00000_00000_00000111110; // lcdwrite 20 62
	HD[2426] = 32'b100111_11011_00000_00000_00000111100; // lcdwrite 27 60
	HD[2427] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2428] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2429] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2430] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2431] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2432] = 32'b100111_10110_00000_00000_00000111110; // lcdwrite 22 62
	HD[2433] = 32'b100111_11001_00000_00000_00000111100; // lcdwrite 25 60
	HD[2434] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2435] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2436] = 32'b000010_10101_00011_0000000000000001; // sw 3 $fp 1
	HD[2437] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2438] = 32'b101000_00000000000000000000100001; // jal sleep
	HD[2439] = 32'b100110_00000000000000000000000000; // lcdclean
	HD[2440] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2441] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2442] = 32'b001111_10110_10111_0000000000000000; // push $ra / menu_opt7_help
	HD[2443] = 32'b100111_00000_00000_00000_00000100000; // lcdwrite 0 32
	HD[2444] = 32'b100111_00001_00000_00000_00001001001; // lcdwrite 1 73
	HD[2445] = 32'b100111_00010_00000_00000_00001101110; // lcdwrite 2 110
	HD[2446] = 32'b100111_00011_00000_00000_00001110011; // lcdwrite 3 115
	HD[2447] = 32'b100111_00100_00000_00000_00001101001; // lcdwrite 4 105
	HD[2448] = 32'b100111_00101_00000_00000_00001110010; // lcdwrite 5 114
	HD[2449] = 32'b100111_00110_00000_00000_00001100001; // lcdwrite 6 97
	HD[2450] = 32'b100111_00111_00000_00000_00000100000; // lcdwrite 7 32
	HD[2451] = 32'b100111_01000_00000_00000_00000101000; // lcdwrite 8 40
	HD[2452] = 32'b100111_01001_00000_00000_00000110001; // lcdwrite 9 49
	HD[2453] = 32'b100111_01010_00000_00000_00000101001; // lcdwrite 10 41
	HD[2454] = 32'b100111_01011_00000_00000_00000100000; // lcdwrite 11 32
	HD[2455] = 32'b100111_01100_00000_00000_00001110000; // lcdwrite 12 112
	HD[2456] = 32'b100111_01101_00000_00000_00001100001; // lcdwrite 13 97
	HD[2457] = 32'b100111_01110_00000_00000_00001110010; // lcdwrite 14 114
	HD[2458] = 32'b100111_01111_00000_00000_00001100001; // lcdwrite 15 97
	HD[2459] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2460] = 32'b100111_10001_00000_00000_00001101001; // lcdwrite 17 105
	HD[2461] = 32'b100111_10010_00000_00000_00001110010; // lcdwrite 18 114
	HD[2462] = 32'b100111_10011_00000_00000_00000100000; // lcdwrite 19 32
	HD[2463] = 32'b100111_10100_00000_00000_00001110000; // lcdwrite 20 112
	HD[2464] = 32'b100111_10101_00000_00000_00001100001; // lcdwrite 21 97
	HD[2465] = 32'b100111_10110_00000_00000_00001110010; // lcdwrite 22 114
	HD[2466] = 32'b100111_10111_00000_00000_00001100001; // lcdwrite 23 97
	HD[2467] = 32'b100111_11000_00000_00000_00000100000; // lcdwrite 24 32
	HD[2468] = 32'b100111_11001_00000_00000_00001101111; // lcdwrite 25 111
	HD[2469] = 32'b100111_11010_00000_00000_00000100000; // lcdwrite 26 32
	HD[2470] = 32'b100111_11011_00000_00000_00001110000; // lcdwrite 27 112
	HD[2471] = 32'b100111_11100_00000_00000_00001110010; // lcdwrite 28 114
	HD[2472] = 32'b100111_11101_00000_00000_00001101111; // lcdwrite 29 111
	HD[2473] = 32'b100111_11110_00000_00000_00001111000; // lcdwrite 30 120
	HD[2474] = 32'b100111_11111_00000_00000_00000101110; // lcdwrite 31 46
	HD[2475] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[2476] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2477] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin17_
	HD[2478] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[2479] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2480] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[2481] = 32'b000111_00010_00000_0000000000000100; // beq 2 $zero _WhileExit17_
	HD[2482] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[2483] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2484] = 32'b001011_00000000000000100110101101; // jump _WhileBegin17_
	HD[2485] = 32'b100111_01001_00000_00000_00000110010; // lcdwrite 9 50 / _WhileExit17_
	HD[2486] = 32'b100111_11011_00000_00000_00001100001; // lcdwrite 27 97
	HD[2487] = 32'b100111_11100_00000_00000_00001101110; // lcdwrite 28 110
	HD[2488] = 32'b100111_11101_00000_00000_00001110100; // lcdwrite 29 116
	HD[2489] = 32'b100111_11110_00000_00000_00000101110; // lcdwrite 30 46
	HD[2490] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2491] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin18_
	HD[2492] = 32'b000101_00000_00011_0000000000000010; // li 3 2
	HD[2493] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2494] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[2495] = 32'b000111_00010_00000_0000000000000100; // beq 2 $zero _WhileExit18_
	HD[2496] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[2497] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2498] = 32'b001011_00000000000000100110111011; // jump _WhileBegin18_
	HD[2499] = 32'b100111_01001_00000_00000_00000110011; // lcdwrite 9 51 / _WhileExit18_
	HD[2500] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2501] = 32'b100111_10001_00000_00000_00001100011; // lcdwrite 17 99
	HD[2502] = 32'b100111_10010_00000_00000_00001101111; // lcdwrite 18 111
	HD[2503] = 32'b100111_10011_00000_00000_00001101110; // lcdwrite 19 110
	HD[2504] = 32'b100111_10100_00000_00000_00001100110; // lcdwrite 20 102
	HD[2505] = 32'b100111_10101_00000_00000_00001101001; // lcdwrite 21 105
	HD[2506] = 32'b100111_10110_00000_00000_00001110010; // lcdwrite 22 114
	HD[2507] = 32'b100111_10111_00000_00000_00001101101; // lcdwrite 23 109
	HD[2508] = 32'b100111_11000_00000_00000_00001100001; // lcdwrite 24 97
	HD[2509] = 32'b100111_11001_00000_00000_00001110010; // lcdwrite 25 114
	HD[2510] = 32'b100111_11010_00000_00000_00000100000; // lcdwrite 26 32
	HD[2511] = 32'b100111_11011_00000_00000_00001101111; // lcdwrite 27 111
	HD[2512] = 32'b100111_11100_00000_00000_00001110000; // lcdwrite 28 112
	HD[2513] = 32'b100111_11101_00000_00000_00001100011; // lcdwrite 29 99
	HD[2514] = 32'b100111_11110_00000_00000_00001100001; // lcdwrite 30 97
	HD[2515] = 32'b100111_11111_00000_00000_00001101111; // lcdwrite 31 111
	HD[2516] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin19_
	HD[2517] = 32'b000101_00000_00011_0000000000000011; // li 3 3
	HD[2518] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2519] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[2520] = 32'b000111_00010_00000_0000000000000100; // beq 2 $zero _WhileExit19_
	HD[2521] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[2522] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2523] = 32'b001011_00000000000000100111010100; // jump _WhileBegin19_
	HD[2524] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _WhileExit19_
	HD[2525] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2526] = 32'b001111_10110_10111_0000000000000000; // push $ra / print_menu
	HD[2527] = 32'b100111_00000_00000_00000_00000100000; // lcdwrite 0 32
	HD[2528] = 32'b100111_00001_00000_00000_00000100000; // lcdwrite 1 32
	HD[2529] = 32'b100111_00010_00000_00000_00001101001; // lcdwrite 2 105
	HD[2530] = 32'b100111_00011_00000_00000_00001101100; // lcdwrite 3 108
	HD[2531] = 32'b100111_00100_00000_00000_00001101111; // lcdwrite 4 111
	HD[2532] = 32'b100111_00101_00000_00000_00001101111; // lcdwrite 5 111
	HD[2533] = 32'b100111_00110_00000_00000_00001110000; // lcdwrite 6 112
	HD[2534] = 32'b100111_00111_00000_00000_00000110011; // lcdwrite 7 51
	HD[2535] = 32'b100111_01000_00000_00000_00000110010; // lcdwrite 8 50
	HD[2536] = 32'b100111_01001_00000_00000_00000100000; // lcdwrite 9 32
	HD[2537] = 32'b100111_01010_00000_00000_00001001101; // lcdwrite 10 77
	HD[2538] = 32'b100111_01011_00000_00000_00001000101; // lcdwrite 11 69
	HD[2539] = 32'b100111_01100_00000_00000_00001001110; // lcdwrite 12 78
	HD[2540] = 32'b100111_01101_00000_00000_00001010101; // lcdwrite 13 85
	HD[2541] = 32'b100111_01110_00000_00000_00000100000; // lcdwrite 14 32
	HD[2542] = 32'b100111_01111_00000_00000_00000100000; // lcdwrite 15 32
	HD[2543] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[2544] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2545] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2546] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin61_
	HD[2547] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2548] = 32'b100111_10001_00000_00000_00001000101; // lcdwrite 17 69
	HD[2549] = 32'b100111_10010_00000_00000_00001111000; // lcdwrite 18 120
	HD[2550] = 32'b100111_10011_00000_00000_00001100101; // lcdwrite 19 101
	HD[2551] = 32'b100111_10100_00000_00000_00001100011; // lcdwrite 20 99
	HD[2552] = 32'b100111_10101_00000_00000_00001110101; // lcdwrite 21 117
	HD[2553] = 32'b100111_10110_00000_00000_00001110100; // lcdwrite 22 116
	HD[2554] = 32'b100111_10111_00000_00000_00001100001; // lcdwrite 23 97
	HD[2555] = 32'b100111_11000_00000_00000_00001110010; // lcdwrite 24 114
	HD[2556] = 32'b100111_11001_00000_00000_00000100000; // lcdwrite 25 32
	HD[2557] = 32'b100111_11010_00000_00000_00001010000; // lcdwrite 26 80
	HD[2558] = 32'b100111_11011_00000_00000_00001110010; // lcdwrite 27 114
	HD[2559] = 32'b100111_11100_00000_00000_00001101111; // lcdwrite 28 111
	HD[2560] = 32'b100111_11101_00000_00000_00001100111; // lcdwrite 29 103
	HD[2561] = 32'b100111_11110_00000_00000_00000101110; // lcdwrite 30 46
	HD[2562] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2563] = 32'b001011_00000000000000101010010010; // jump _IfExit61_
	HD[2564] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin61_
	HD[2565] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[2566] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2567] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin62_
	HD[2568] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2569] = 32'b100111_10001_00000_00000_00001000101; // lcdwrite 17 69
	HD[2570] = 32'b100111_10010_00000_00000_00001110011; // lcdwrite 18 115
	HD[2571] = 32'b100111_10011_00000_00000_00001100011; // lcdwrite 19 99
	HD[2572] = 32'b100111_10100_00000_00000_00001110010; // lcdwrite 20 114
	HD[2573] = 32'b100111_10101_00000_00000_00001100101; // lcdwrite 21 101
	HD[2574] = 32'b100111_10110_00000_00000_00001110110; // lcdwrite 22 118
	HD[2575] = 32'b100111_10111_00000_00000_00001100101; // lcdwrite 23 101
	HD[2576] = 32'b100111_11000_00000_00000_00001110010; // lcdwrite 24 114
	HD[2577] = 32'b100111_11001_00000_00000_00000100000; // lcdwrite 25 32
	HD[2578] = 32'b100111_11010_00000_00000_00001010000; // lcdwrite 26 80
	HD[2579] = 32'b100111_11011_00000_00000_00001110010; // lcdwrite 27 114
	HD[2580] = 32'b100111_11100_00000_00000_00001101111; // lcdwrite 28 111
	HD[2581] = 32'b100111_11101_00000_00000_00001100111; // lcdwrite 29 103
	HD[2582] = 32'b100111_11110_00000_00000_00000101110; // lcdwrite 30 46
	HD[2583] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2584] = 32'b001011_00000000000000101010010010; // jump _IfExit62_
	HD[2585] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin62_
	HD[2586] = 32'b000101_00000_00011_0000000000000010; // li 3 2
	HD[2587] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2588] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin63_
	HD[2589] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2590] = 32'b100111_10001_00000_00000_00001010010; // lcdwrite 17 82
	HD[2591] = 32'b100111_10010_00000_00000_00001100101; // lcdwrite 18 101
	HD[2592] = 32'b100111_10011_00000_00000_00001101110; // lcdwrite 19 110
	HD[2593] = 32'b100111_10100_00000_00000_00001101111; // lcdwrite 20 111
	HD[2594] = 32'b100111_10101_00000_00000_00001101101; // lcdwrite 21 109
	HD[2595] = 32'b100111_10110_00000_00000_00001100101; // lcdwrite 22 101
	HD[2596] = 32'b100111_10111_00000_00000_00001100001; // lcdwrite 23 97
	HD[2597] = 32'b100111_11000_00000_00000_00001110010; // lcdwrite 24 114
	HD[2598] = 32'b100111_11001_00000_00000_00000100000; // lcdwrite 25 32
	HD[2599] = 32'b100111_11010_00000_00000_00001010000; // lcdwrite 26 80
	HD[2600] = 32'b100111_11011_00000_00000_00001110010; // lcdwrite 27 114
	HD[2601] = 32'b100111_11100_00000_00000_00001101111; // lcdwrite 28 111
	HD[2602] = 32'b100111_11101_00000_00000_00001100111; // lcdwrite 29 103
	HD[2603] = 32'b100111_11110_00000_00000_00000101110; // lcdwrite 30 46
	HD[2604] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2605] = 32'b001011_00000000000000101010010010; // jump _IfExit63_
	HD[2606] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin63_
	HD[2607] = 32'b000101_00000_00011_0000000000000011; // li 3 3
	HD[2608] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2609] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin64_
	HD[2610] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2611] = 32'b100111_10001_00000_00000_00001000100; // lcdwrite 17 68
	HD[2612] = 32'b100111_10010_00000_00000_00001100101; // lcdwrite 18 101
	HD[2613] = 32'b100111_10011_00000_00000_00001101100; // lcdwrite 19 108
	HD[2614] = 32'b100111_10100_00000_00000_00001100101; // lcdwrite 20 101
	HD[2615] = 32'b100111_10101_00000_00000_00001110100; // lcdwrite 21 116
	HD[2616] = 32'b100111_10110_00000_00000_00001100001; // lcdwrite 22 97
	HD[2617] = 32'b100111_10111_00000_00000_00001110010; // lcdwrite 23 114
	HD[2618] = 32'b100111_11000_00000_00000_00000100000; // lcdwrite 24 32
	HD[2619] = 32'b100111_11001_00000_00000_00000100000; // lcdwrite 25 32
	HD[2620] = 32'b100111_11010_00000_00000_00001010000; // lcdwrite 26 80
	HD[2621] = 32'b100111_11011_00000_00000_00001110010; // lcdwrite 27 114
	HD[2622] = 32'b100111_11100_00000_00000_00001101111; // lcdwrite 28 111
	HD[2623] = 32'b100111_11101_00000_00000_00001100111; // lcdwrite 29 103
	HD[2624] = 32'b100111_11110_00000_00000_00000101110; // lcdwrite 30 46
	HD[2625] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2626] = 32'b001011_00000000000000101010010010; // jump _IfExit64_
	HD[2627] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin64_
	HD[2628] = 32'b000101_00000_00011_0000000000000100; // li 3 4
	HD[2629] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2630] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin65_
	HD[2631] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2632] = 32'b100111_10001_00000_00000_00001001100; // lcdwrite 17 76
	HD[2633] = 32'b100111_10010_00000_00000_00001101001; // lcdwrite 18 105
	HD[2634] = 32'b100111_10011_00000_00000_00001110011; // lcdwrite 19 115
	HD[2635] = 32'b100111_10100_00000_00000_00001110100; // lcdwrite 20 116
	HD[2636] = 32'b100111_10101_00000_00000_00001100001; // lcdwrite 21 97
	HD[2637] = 32'b100111_10110_00000_00000_00001110010; // lcdwrite 22 114
	HD[2638] = 32'b100111_10111_00000_00000_00000100000; // lcdwrite 23 32
	HD[2639] = 32'b100111_11000_00000_00000_00000100000; // lcdwrite 24 32
	HD[2640] = 32'b100111_11001_00000_00000_00000100000; // lcdwrite 25 32
	HD[2641] = 32'b100111_11010_00000_00000_00001010000; // lcdwrite 26 80
	HD[2642] = 32'b100111_11011_00000_00000_00001110010; // lcdwrite 27 114
	HD[2643] = 32'b100111_11100_00000_00000_00001101111; // lcdwrite 28 111
	HD[2644] = 32'b100111_11101_00000_00000_00001100111; // lcdwrite 29 103
	HD[2645] = 32'b100111_11110_00000_00000_00000101110; // lcdwrite 30 46
	HD[2646] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2647] = 32'b001011_00000000000000101010010010; // jump _IfExit65_
	HD[2648] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin65_
	HD[2649] = 32'b000101_00000_00011_0000000000000101; // li 3 5
	HD[2650] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2651] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin66_
	HD[2652] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2653] = 32'b100111_10001_00000_00000_00001010010; // lcdwrite 17 82
	HD[2654] = 32'b100111_10010_00000_00000_00001100101; // lcdwrite 18 101
	HD[2655] = 32'b100111_10011_00000_00000_00001101001; // lcdwrite 19 105
	HD[2656] = 32'b100111_10100_00000_00000_00001101110; // lcdwrite 20 110
	HD[2657] = 32'b100111_10101_00000_00000_00001101001; // lcdwrite 21 105
	HD[2658] = 32'b100111_10110_00000_00000_00001100011; // lcdwrite 22 99
	HD[2659] = 32'b100111_10111_00000_00000_00001101001; // lcdwrite 23 105
	HD[2660] = 32'b100111_11000_00000_00000_00001100001; // lcdwrite 24 97
	HD[2661] = 32'b100111_11001_00000_00000_00001110010; // lcdwrite 25 114
	HD[2662] = 32'b100111_11010_00000_00000_00000100000; // lcdwrite 26 32
	HD[2663] = 32'b100111_11011_00000_00000_00001010011; // lcdwrite 27 83
	HD[2664] = 32'b100111_11100_00000_00000_00000101110; // lcdwrite 28 46
	HD[2665] = 32'b100111_11101_00000_00000_00001001111; // lcdwrite 29 79
	HD[2666] = 32'b100111_11110_00000_00000_00000101110; // lcdwrite 30 46
	HD[2667] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2668] = 32'b001011_00000000000000101010010010; // jump _IfExit66_
	HD[2669] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin66_
	HD[2670] = 32'b000101_00000_00011_0000000000000110; // li 3 6
	HD[2671] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2672] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin67_
	HD[2673] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32
	HD[2674] = 32'b100111_10001_00000_00000_00001000100; // lcdwrite 17 68
	HD[2675] = 32'b100111_10010_00000_00000_00001100101; // lcdwrite 18 101
	HD[2676] = 32'b100111_10011_00000_00000_00001110011; // lcdwrite 19 115
	HD[2677] = 32'b100111_10100_00000_00000_00001101100; // lcdwrite 20 108
	HD[2678] = 32'b100111_10101_00000_00000_00001101001; // lcdwrite 21 105
	HD[2679] = 32'b100111_10110_00000_00000_00001100111; // lcdwrite 22 103
	HD[2680] = 32'b100111_10111_00000_00000_00001100001; // lcdwrite 23 97
	HD[2681] = 32'b100111_11000_00000_00000_00001110010; // lcdwrite 24 114
	HD[2682] = 32'b100111_11001_00000_00000_00000100000; // lcdwrite 25 32
	HD[2683] = 32'b100111_11010_00000_00000_00000100000; // lcdwrite 26 32
	HD[2684] = 32'b100111_11011_00000_00000_00001010011; // lcdwrite 27 83
	HD[2685] = 32'b100111_11100_00000_00000_00000101110; // lcdwrite 28 46
	HD[2686] = 32'b100111_11101_00000_00000_00001001111; // lcdwrite 29 79
	HD[2687] = 32'b100111_11110_00000_00000_00000101110; // lcdwrite 30 46
	HD[2688] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2689] = 32'b001011_00000000000000101010010010; // jump _IfExit67_
	HD[2690] = 32'b100111_10000_00000_00000_00000100000; // lcdwrite 16 32 / _ElseBegin67_
	HD[2691] = 32'b100111_10001_00000_00000_00000101101; // lcdwrite 17 45
	HD[2692] = 32'b100111_10010_00000_00000_00000101101; // lcdwrite 18 45
	HD[2693] = 32'b100111_10011_00000_00000_00001000010; // lcdwrite 19 66
	HD[2694] = 32'b100111_10100_00000_00000_00001100001; // lcdwrite 20 97
	HD[2695] = 32'b100111_10101_00000_00000_00001110011; // lcdwrite 21 115
	HD[2696] = 32'b100111_10110_00000_00000_00001101000; // lcdwrite 22 104
	HD[2697] = 32'b100111_10111_00000_00000_00000100000; // lcdwrite 23 32
	HD[2698] = 32'b100111_11000_00000_00000_00000100000; // lcdwrite 24 32
	HD[2699] = 32'b100111_11001_00000_00000_00001001000; // lcdwrite 25 72
	HD[2700] = 32'b100111_11010_00000_00000_00001100101; // lcdwrite 26 101
	HD[2701] = 32'b100111_11011_00000_00000_00001101100; // lcdwrite 27 108
	HD[2702] = 32'b100111_11100_00000_00000_00001110000; // lcdwrite 28 112
	HD[2703] = 32'b100111_11101_00000_00000_00000101101; // lcdwrite 29 45
	HD[2704] = 32'b100111_11110_00000_00000_00000101101; // lcdwrite 30 45
	HD[2705] = 32'b100111_11111_00000_00000_00000100000; // lcdwrite 31 32
	HD[2706] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _IfExit67_ _IfExit66_ _IfExit65_ _IfExit64_ _IfExit63_ _IfExit62_ _IfExit61_
	HD[2707] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2708] = 32'b001111_10110_10111_0000000000000000; // push $ra / tela_prox
	HD[2709] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2710] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[2711] = 32'b000101_00000_00010_0000000000000111; // li 2 7
	HD[2712] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[2713] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[2714] = 32'b000001_10101_00011_0000000000000010; // lw 3 $fp 2
	HD[2715] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2716] = 32'b000111_00010_00000_0000000000000110; // beq 2 $zero _ElseBegin68_
	HD[2717] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[2718] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[2719] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2720] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2721] = 32'b001011_00000000000000101010100111; // jump _IfExit68_
	HD[2722] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin68_
	HD[2723] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[2724] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[2725] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2726] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2727] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _IfExit68_
	HD[2728] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2729] = 32'b001111_10110_10111_0000000000000000; // push $ra / tela_ant
	HD[2730] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2731] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[2732] = 32'b000101_00000_00010_0000000000000111; // li 2 7
	HD[2733] = 32'b000010_10101_00010_0000000000000010; // sw 2 $fp 2
	HD[2734] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[2735] = 32'b000001_10101_00011_0000000000000001; // lw 3 $fp 1
	HD[2736] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2737] = 32'b000111_00010_00000_0000000000000110; // beq 2 $zero _ElseBegin69_
	HD[2738] = 32'b000001_10101_00010_0000000000000010; // lw 2 $fp 2
	HD[2739] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[2740] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2741] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2742] = 32'b001011_00000000000000101010111100; // jump _IfExit69_
	HD[2743] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin69_
	HD[2744] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[2745] = 32'b000000_00010_10100_00000_00000_010000; // move $rv 2
	HD[2746] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2747] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2748] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _IfExit69_
	HD[2749] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2750] = 32'b001111_10110_10111_0000000000000000; // push $ra / bash_OS
	HD[2751] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2752] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2753] = 32'b000101_00000_00010_0000000000000001; // li 2 1 / _WhileBegin20_
	HD[2754] = 32'b000111_00010_00000_0000000001100010; // beq 2 $zero _WhileExit20_
	HD[2755] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[2756] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2757] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2758] = 32'b101000_00000000000000100111011110; // jal print_menu
	HD[2759] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2760] = 32'b001001_00000_00010_0000000000000000; // in 2
	HD[2761] = 32'b000010_10101_00010_0000000000000001; // sw 2 $fp 1
	HD[2762] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1
	HD[2763] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[2764] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2765] = 32'b000111_00010_00000_0000000000001001; // beq 2 $zero _ElseBegin70_
	HD[2766] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[2767] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2768] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2769] = 32'b101000_00000000000000101010010100; // jal tela_prox
	HD[2770] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2771] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[2772] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2773] = 32'b001011_00000000000000101100100011; // jump _IfExit70_
	HD[2774] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _ElseBegin70_
	HD[2775] = 32'b000101_00000_00011_0000000000000010; // li 3 2
	HD[2776] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2777] = 32'b000111_00010_00000_0000000000001001; // beq 2 $zero _ElseBegin71_
	HD[2778] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[2779] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2780] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2781] = 32'b101000_00000000000000101010101001; // jal tela_ant
	HD[2782] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2783] = 32'b000000_10100_00010_00000_00000_010000; // move 2 $rv
	HD[2784] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2785] = 32'b001011_00000000000000101100100011; // jump _IfExit71_
	HD[2786] = 32'b000001_10101_00010_0000000000000001; // lw 2 $fp 1 / _ElseBegin71_
	HD[2787] = 32'b000101_00000_00011_0000000000000011; // li 3 3
	HD[2788] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2789] = 32'b000111_00010_00000_0000000000111110; // beq 2 $zero _IfExit72_
	HD[2790] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[2791] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[2792] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2793] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin73_
	HD[2794] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2795] = 32'b101000_00000000000000010111111101; // jal menu_opt0_executar_prog
	HD[2796] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2797] = 32'b001011_00000000000000101100100011; // jump _IfExit73_
	HD[2798] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin73_
	HD[2799] = 32'b000101_00000_00011_0000000000000001; // li 3 1
	HD[2800] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2801] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin74_
	HD[2802] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2803] = 32'b101000_00000000000000011010001010; // jal menu_opt1_escrever_prog
	HD[2804] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2805] = 32'b001011_00000000000000101100100011; // jump _IfExit74_
	HD[2806] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin74_
	HD[2807] = 32'b000101_00000_00011_0000000000000010; // li 3 2
	HD[2808] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2809] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin75_
	HD[2810] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2811] = 32'b101000_00000000000000011101101001; // jal menu_opt2_renomear_prog
	HD[2812] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2813] = 32'b001011_00000000000000101100100011; // jump _IfExit75_
	HD[2814] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin75_
	HD[2815] = 32'b000101_00000_00011_0000000000000011; // li 3 3
	HD[2816] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2817] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin76_
	HD[2818] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2819] = 32'b101000_00000000000000100001000110; // jal menu_opt3_deletar_prog
	HD[2820] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2821] = 32'b001011_00000000000000101100100011; // jump _IfExit76_
	HD[2822] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin76_
	HD[2823] = 32'b000101_00000_00011_0000000000000100; // li 3 4
	HD[2824] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2825] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin77_
	HD[2826] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2827] = 32'b101000_00000000000000100010111111; // jal menu_opt4_listar_prog
	HD[2828] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2829] = 32'b001011_00000000000000101100100011; // jump _IfExit77_
	HD[2830] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin77_
	HD[2831] = 32'b000101_00000_00011_0000000000000101; // li 3 5
	HD[2832] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2833] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin78_
	HD[2834] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2835] = 32'b101000_00000000000000100100100011; // jal menu_opt5_reiniciar
	HD[2836] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2837] = 32'b001011_00000000000000101100100011; // jump _IfExit78_
	HD[2838] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin78_
	HD[2839] = 32'b000101_00000_00011_0000000000000110; // li 3 6
	HD[2840] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
	HD[2841] = 32'b000111_00010_00000_0000000000000111; // beq 2 $zero _ElseBegin79_
	HD[2842] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2
	HD[2843] = 32'b101000_00000000000000100101011010; // jal menu_opt6_desligar
	HD[2844] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2845] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2846] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2847] = 32'b001011_00000000000000101100100011; // jump _IfExit79_
	HD[2848] = 32'b000011_10101_10101_0000000000000010; // addi $fp $fp 2 / _ElseBegin79_
	HD[2849] = 32'b101000_00000000000000100110001010; // jal menu_opt7_help
	HD[2850] = 32'b000100_10101_10101_0000000000000010; // subi $fp $fp 2
	HD[2851] = 32'b001011_00000000000000101011000001; // jump _WhileBegin20_ / _IfExit79_ _IfExit78_ _IfExit77_ _IfExit76_ _IfExit75_ _IfExit74_ _IfExit73_ _IfExit72_ _IfExit71_ _IfExit70_
	HD[2852] = 32'b010000_10110_10111_0000000000000000; // pop $ra / _WhileExit20_
	HD[2853] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2854] = 32'b001111_10110_10111_0000000000000000; // push $ra / init_global
	HD[2855] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2856] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2857] = 32'b000101_00000_00010_0000000000001111; // li 2 15
	HD[2858] = 32'b000010_00000_00010_0000000000000000; // sw 2 $global 0
	HD[2859] = 32'b000101_00000_00010_0000101110111000; // li 2 3000
	HD[2860] = 32'b000010_00000_00010_0000000000000001; // sw 2 $global 1
	HD[2861] = 32'b000101_00000_00010_0000000100000000; // li 2 256
	HD[2862] = 32'b000010_00000_00010_0000000000000010; // sw 2 $global 2
	HD[2863] = 32'b000101_00000_00010_0000100000000000; // li 2 2048
	HD[2864] = 32'b000010_00000_00010_0000000000000011; // sw 2 $global 3
	HD[2865] = 32'b000101_00000_00010_0000000100000000; // li 2 256
	HD[2866] = 32'b000010_00000_00010_0000000000000100; // sw 2 $global 4
	HD[2867] = 32'b000101_00000_00010_0000000000100000; // li 2 32
	HD[2868] = 32'b000010_00000_00010_0000000000000101; // sw 2 $global 5
	HD[2869] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2870] = 32'b000010_00000_00010_0000000000000110; // sw 2 $global 6
	HD[2871] = 32'b000101_00000_00010_0000000000001010; // li 2 10
	HD[2872] = 32'b000010_00000_00010_0000000000000111; // sw 2 $global 7
	HD[2873] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2874] = 32'b000010_00000_00010_0000000000001000; // sw 2 $global 8
	HD[2875] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin21_
	HD[2876] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[2877] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[2878] = 32'b000111_00010_00000_0000000000001001; // beq 2 $zero _WhileExit21_
	HD[2879] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2880] = 32'b000001_10101_00011_0000000000000000; // lw 3 $fp 0
	HD[2881] = 32'b000000_00011_00000_00011_00000_000101; // add 3 3 $global
	HD[2882] = 32'b000010_00011_00010_0000000000001001; // sw 2 3 9
	HD[2883] = 32'b000001_10101_00010_0000000000000000; // lw 2 $fp 0
	HD[2884] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[2885] = 32'b000010_10101_00010_0000000000000000; // sw 2 $fp 0
	HD[2886] = 32'b001011_00000000000000101100111011; // jump _WhileBegin21_
	HD[2887] = 32'b000101_00000_00010_0000000000000000; // li 2 0 / _WhileExit21_
	HD[2888] = 32'b000010_00000_00010_0000000000010011; // sw 2 $global 19
	HD[2889] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2890] = 32'b000010_00000_00010_0000000000010100; // sw 2 $global 20
	HD[2891] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2892] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[2893] = 32'b000010_00000_00010_0000000000010101; // sw 2 $global 21
	HD[2894] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2895] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[2896] = 32'b000010_00000_00010_0000000000010110; // sw 2 $global 22
	HD[2897] = 32'b000101_00000_00010_0000000000000011; // li 2 3
	HD[2898] = 32'b000010_00000_00010_0000000000010111; // sw 2 $global 23
	HD[2899] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2900] = 32'b000010_00000_00010_0000000000011000; // sw 2 $global 24
	HD[2901] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2902] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
	HD[2903] = 32'b000010_00000_00010_0000000000011001; // sw 2 $global 25
	HD[2904] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2905] = 32'b000100_00010_00010_0000000000000010; // subi 2 2 2
	HD[2906] = 32'b000010_00000_00010_0000000000011010; // sw 2 $global 26
	HD[2907] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2908] = 32'b000100_00010_00010_0000000000000011; // subi 2 2 3
	HD[2909] = 32'b000010_00000_00010_0000000000011011; // sw 2 $global 27
	HD[2910] = 32'b000101_00000_00010_0000000000000011; // li 2 3
	HD[2911] = 32'b000010_00000_00010_0000000000011100; // sw 2 $global 28
	HD[2912] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[2913] = 32'b000010_00000_00010_0000000000011101; // sw 2 $global 29
	HD[2914] = 32'b000101_00000_00010_0000000000000001; // li 2 1
	HD[2915] = 32'b000010_00000_00010_0000000000011110; // sw 2 $global 30
	HD[2916] = 32'b000101_00000_00010_0000000000000010; // li 2 2
	HD[2917] = 32'b000010_00000_00010_0000000000011111; // sw 2 $global 31
	HD[2918] = 32'b000101_00000_00010_0000000000000011; // li 2 3
	HD[2919] = 32'b000010_00000_00010_0000000000100000; // sw 2 $global 32
	HD[2920] = 32'b010000_10110_10111_0000000000000000; // pop $ra
	HD[2921] = 32'b000000_10111_00000_00000_00000_010100; // jr $ra
	HD[2922] = 32'b101000_00000000000000101100100110; // jal init_global / main
	HD[2923] = 32'b101000_00000000000000101010111110; // jal bash_OS
	HD[2924] = 32'b11111111111111111111111111111111; // halt / _halt_
	
	
	/* Programa 01 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 3075> */
	HD[3075] = 32'b000011_11011_11101_0000000000001010; // addi $fp $global 10
	HD[3076] = 32'b001011_00000000000000110000110010; // jump main
	HD[3077] = 32'b001111_11110_11111_0000000000000000; // push $ra / minloc
	HD[3078] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1
	HD[3079] = 32'b000010_11101_01010_0000000000000101; // sw 10 $fp 5
	HD[3080] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[3081] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[3082] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[3083] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[3084] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[3085] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1
	HD[3086] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[3087] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[3088] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _WhileBegin0_
	HD[3089] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[3090] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[3091] = 32'b000111_01010_00000_0000000000010011; // beq 10 $zero _WhileExit0_
	HD[3092] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[3093] = 32'b000001_11101_01011_0000000000000011; // lw 11 $fp 3
	HD[3094] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[3095] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[3096] = 32'b000001_11101_01011_0000000000000100; // lw 11 $fp 4
	HD[3097] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[3098] = 32'b000111_01010_00000_0000000000001000; // beq 10 $zero _IfExit0_
	HD[3099] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[3100] = 32'b000001_11101_01011_0000000000000011; // lw 11 $fp 3
	HD[3101] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[3102] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[3103] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[3104] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3
	HD[3105] = 32'b000010_11101_01010_0000000000000101; // sw 10 $fp 5
	HD[3106] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _IfExit0_
	HD[3107] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[3108] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[3109] = 32'b001011_00000000000000101111000101; // jump _WhileBegin0_
	HD[3110] = 32'b000001_11101_01010_0000000000000101; // lw 10 $fp 5 / _WhileExit0_
	HD[3111] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[3112] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[3113] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[3114] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[3115] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[3116] = 32'b001111_11110_11111_0000000000000000; // push $ra / sort
	HD[3117] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1
	HD[3118] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[3119] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _WhileBegin1_
	HD[3120] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[3121] = 32'b000100_01011_01011_0000000000000001; // subi 11 11 1
	HD[3122] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[3123] = 32'b000111_01010_00000_0000000000100010; // beq 10 $zero _WhileExit1_
	HD[3124] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[3125] = 32'b000001_11101_01011_0000000000000011; // lw 11 $fp 3
	HD[3126] = 32'b000001_11101_01100_0000000000000010; // lw 12 $fp 2
	HD[3127] = 32'b000011_11101_11101_0000000000000110; // addi $fp $fp 6
	HD[3128] = 32'b000010_11101_01100_0000000000000010; // sw 12 $fp 2
	HD[3129] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[3130] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[3131] = 32'b001100_00000000000000101110111010; // jal minloc
	HD[3132] = 32'b000100_11101_11101_0000000000000110; // subi $fp $fp 6
	HD[3133] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[3134] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[3135] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[3136] = 32'b000001_11101_01011_0000000000000100; // lw 11 $fp 4
	HD[3137] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[3138] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[3139] = 32'b000010_11101_01010_0000000000000101; // sw 10 $fp 5
	HD[3140] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[3141] = 32'b000001_11101_01011_0000000000000011; // lw 11 $fp 3
	HD[3142] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[3143] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[3144] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[3145] = 32'b000001_11101_01100_0000000000000100; // lw 12 $fp 4
	HD[3146] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[3147] = 32'b000010_01011_01010_0000000000000000; // sw 10 11 0
	HD[3148] = 32'b000001_11101_01010_0000000000000101; // lw 10 $fp 5
	HD[3149] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[3150] = 32'b000001_11101_01100_0000000000000011; // lw 12 $fp 3
	HD[3151] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[3152] = 32'b000010_01011_01010_0000000000000000; // sw 10 11 0
	HD[3153] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3
	HD[3154] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[3155] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[3156] = 32'b001011_00000000000000101111100100; // jump _WhileBegin1_
	HD[3157] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit1_
	HD[3158] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[3159] = 32'b001111_11110_11111_0000000000000000; // push $ra / inputVector
	HD[3160] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[3161] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[3162] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin2_
	HD[3163] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[3164] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[3165] = 32'b000111_01010_00000_0000000000001011; // beq 10 $zero _WhileExit2_
	HD[3166] = 32'b101101_00000000000000000000000100; // syscall 0
	HD[3167] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[3168] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[3169] = 32'b000001_11101_01100_0000000000000010; // lw 12 $fp 2
	HD[3170] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[3171] = 32'b000010_01011_01010_0000000000000000; // sw 10 11 0
	HD[3172] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[3173] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[3174] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[3175] = 32'b001011_00000000000000110000001111; // jump _WhileBegin2_
	HD[3176] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit2_
	HD[3177] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[3178] = 32'b001111_11110_11111_0000000000000000; // push $ra / outputVector
	HD[3179] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[3180] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[3181] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin3_
	HD[3182] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[3183] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[3184] = 32'b000111_01010_00000_0000000000001011; // beq 10 $zero _WhileExit3_
	HD[3185] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[3186] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[3187] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[3188] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[3189] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[3190] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[3191] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[3192] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[3193] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[3194] = 32'b001011_00000000000000110000100010; // jump _WhileBegin3_
	HD[3195] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit3_
	HD[3196] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[3197] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0 / main
	HD[3198] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[3199] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[3200] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[3201] = 32'b001100_00000000000000110000001100; // jal inputVector
	HD[3202] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0
	HD[3203] = 32'b000101_00000_01011_0000000000000000; // li 11 0
	HD[3204] = 32'b000101_00000_01100_0000000000001010; // li 12 10
	HD[3205] = 32'b000010_11101_01100_0000000000000010; // sw 12 $fp 2
	HD[3206] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[3207] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[3208] = 32'b001100_00000000000000101111100001; // jal sort
	HD[3209] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0
	HD[3210] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[3211] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[3212] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[3213] = 32'b001100_00000000000000110000011111; // jal outputVector
	HD[3214] = 32'b101100_00000000000000000000001111; // return / _halt_

	/* Programa 02 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 4099> */
	HD[4099] = 32'b000011_11011_11101_0000000000001010; // addi $fp $global 10
	HD[4100] = 32'b001011_00000000000000110010001011; // jump main
	HD[4101] = 32'b001111_11110_11111_0000000000000000; // push $ra / minloc
	HD[4102] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1
	HD[4103] = 32'b000010_11101_01010_0000000000000101; // sw 10 $fp 5
	HD[4104] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[4105] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[4106] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[4107] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[4108] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[4109] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1
	HD[4110] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[4111] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[4112] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _WhileBegin0_
	HD[4113] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[4114] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[4115] = 32'b000111_01010_00000_0000000000010011; // beq 10 $zero _WhileExit0_
	HD[4116] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[4117] = 32'b000001_11101_01011_0000000000000011; // lw 11 $fp 3
	HD[4118] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[4119] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[4120] = 32'b000001_11101_01011_0000000000000100; // lw 11 $fp 4
	HD[4121] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[4122] = 32'b000111_01010_00000_0000000000001000; // beq 10 $zero _IfExit0_
	HD[4123] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[4124] = 32'b000001_11101_01011_0000000000000011; // lw 11 $fp 3
	HD[4125] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[4126] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[4127] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[4128] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3
	HD[4129] = 32'b000010_11101_01010_0000000000000101; // sw 10 $fp 5
	HD[4130] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _IfExit0_
	HD[4131] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[4132] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[4133] = 32'b001011_00000000000000101111000101; // jump _WhileBegin0_
	HD[4134] = 32'b000001_11101_01010_0000000000000101; // lw 10 $fp 5 / _WhileExit0_
	HD[4135] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[4136] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[4137] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4138] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[4139] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4140] = 32'b001111_11110_11111_0000000000000000; // push $ra / sort
	HD[4141] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1
	HD[4142] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[4143] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _WhileBegin1_
	HD[4144] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[4145] = 32'b000100_01011_01011_0000000000000001; // subi 11 11 1
	HD[4146] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[4147] = 32'b000111_01010_00000_0000000000100010; // beq 10 $zero _WhileExit1_
	HD[4148] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[4149] = 32'b000001_11101_01011_0000000000000011; // lw 11 $fp 3
	HD[4150] = 32'b000001_11101_01100_0000000000000010; // lw 12 $fp 2
	HD[4151] = 32'b000011_11101_11101_0000000000000110; // addi $fp $fp 6
	HD[4152] = 32'b000010_11101_01100_0000000000000010; // sw 12 $fp 2
	HD[4153] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[4154] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[4155] = 32'b001100_00000000000000101110111010; // jal minloc
	HD[4156] = 32'b000100_11101_11101_0000000000000110; // subi $fp $fp 6
	HD[4157] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[4158] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[4159] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[4160] = 32'b000001_11101_01011_0000000000000100; // lw 11 $fp 4
	HD[4161] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[4162] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[4163] = 32'b000010_11101_01010_0000000000000101; // sw 10 $fp 5
	HD[4164] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[4165] = 32'b000001_11101_01011_0000000000000011; // lw 11 $fp 3
	HD[4166] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[4167] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[4168] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[4169] = 32'b000001_11101_01100_0000000000000100; // lw 12 $fp 4
	HD[4170] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[4171] = 32'b000010_01011_01010_0000000000000000; // sw 10 11 0
	HD[4172] = 32'b000001_11101_01010_0000000000000101; // lw 10 $fp 5
	HD[4173] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[4174] = 32'b000001_11101_01100_0000000000000011; // lw 12 $fp 3
	HD[4175] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[4176] = 32'b000010_01011_01010_0000000000000000; // sw 10 11 0
	HD[4177] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3
	HD[4178] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[4179] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[4180] = 32'b001011_00000000000000101111100100; // jump _WhileBegin1_
	HD[4181] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit1_
	HD[4182] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4183] = 32'b001111_11110_11111_0000000000000000; // push $ra / buscaBinariaInterno
	HD[4184] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[4185] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[4186] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[4187] = 32'b000101_00000_01011_0000000000000010; // li 11 2
	HD[4188] = 32'b000000_01010_01011_01010_00000_001000; // div 10 10 11
	HD[4189] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[4190] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[4191] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[4192] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[4193] = 32'b000111_01010_00000_0000000000000101; // beq 10 $zero _ElseBegin1_
	HD[4194] = 32'b000101_00000_11100_0000000000000000; // li $rv 0
	HD[4195] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[4196] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4197] = 32'b001011_00000000000000110001010001; // jump _IfExit1_
	HD[4198] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _ElseBegin1_
	HD[4199] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[4200] = 32'b000001_11101_01100_0000000000000100; // lw 12 $fp 4
	HD[4201] = 32'b000100_01100_01100_0000000000000001; // subi 12 12 1
	HD[4202] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[4203] = 32'b000001_01011_01011_0000000000000000; // lw 11 11 0
	HD[4204] = 32'b000000_01010_01011_01010_00000_010010; // sgt 10 10 11
	HD[4205] = 32'b000111_01010_00000_0000000000010010; // beq 10 $zero _ElseBegin2_
	HD[4206] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[4207] = 32'b000001_11101_01011_0000000000000100; // lw 11 $fp 4
	HD[4208] = 32'b000011_01011_01011_0000000000000001; // addi 11 11 1
	HD[4209] = 32'b000001_11101_01100_0000000000000010; // lw 12 $fp 2
	HD[4210] = 32'b000001_11101_01101_0000000000000011; // lw 13 $fp 3
	HD[4211] = 32'b000011_11101_11101_0000000000000101; // addi $fp $fp 5
	HD[4212] = 32'b000010_11101_01101_0000000000000011; // sw 13 $fp 3
	HD[4213] = 32'b000010_11101_01100_0000000000000010; // sw 12 $fp 2
	HD[4214] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[4215] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[4216] = 32'b001100_00000000000000110000001100; // jal buscaBinariaInterno
	HD[4217] = 32'b000100_11101_11101_0000000000000101; // subi $fp $fp 5
	HD[4218] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[4219] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[4220] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[4221] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4222] = 32'b001011_00000000000000110001010001; // jump _IfExit2_
	HD[4223] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _ElseBegin2_
	HD[4224] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[4225] = 32'b000001_11101_01100_0000000000000100; // lw 12 $fp 4
	HD[4226] = 32'b000100_01100_01100_0000000000000001; // subi 12 12 1
	HD[4227] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[4228] = 32'b000001_01011_01011_0000000000000000; // lw 11 11 0
	HD[4229] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[4230] = 32'b000111_01010_00000_0000000000010010; // beq 10 $zero _ElseBegin3_
	HD[4231] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[4232] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[4233] = 32'b000001_11101_01100_0000000000000100; // lw 12 $fp 4
	HD[4234] = 32'b000100_01100_01100_0000000000000001; // subi 12 12 1
	HD[4235] = 32'b000001_11101_01101_0000000000000011; // lw 13 $fp 3
	HD[4236] = 32'b000011_11101_11101_0000000000000101; // addi $fp $fp 5
	HD[4237] = 32'b000010_11101_01101_0000000000000011; // sw 13 $fp 3
	HD[4238] = 32'b000010_11101_01100_0000000000000010; // sw 12 $fp 2
	HD[4239] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[4240] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[4241] = 32'b001100_00000000000000110000001100; // jal buscaBinariaInterno
	HD[4242] = 32'b000100_11101_11101_0000000000000101; // subi $fp $fp 5
	HD[4243] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[4244] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[4245] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[4246] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4247] = 32'b001011_00000000000000110001010001; // jump _IfExit3_
	HD[4248] = 32'b000001_11101_01010_0000000000000100; // lw 10 $fp 4 / _ElseBegin3_
	HD[4249] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[4250] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[4251] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4252] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit3_ _IfExit2_ _IfExit1_
	HD[4253] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4254] = 32'b001111_11110_11111_0000000000000000; // push $ra / buscaBinaria
	HD[4255] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[4256] = 32'b000101_00000_01011_0000000000000001; // li 11 1
	HD[4257] = 32'b000001_11101_01100_0000000000000001; // lw 12 $fp 1
	HD[4258] = 32'b000001_11101_01101_0000000000000010; // lw 13 $fp 2
	HD[4259] = 32'b000011_11101_11101_0000000000000011; // addi $fp $fp 3
	HD[4260] = 32'b000010_11101_01101_0000000000000011; // sw 13 $fp 3
	HD[4261] = 32'b000010_11101_01100_0000000000000010; // sw 12 $fp 2
	HD[4262] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[4263] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[4264] = 32'b001100_00000000000000110000001100; // jal buscaBinariaInterno
	HD[4265] = 32'b000100_11101_11101_0000000000000011; // subi $fp $fp 3
	HD[4266] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[4267] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[4268] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[4269] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4270] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[4271] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4272] = 32'b001111_11110_11111_0000000000000000; // push $ra / inputVector
	HD[4273] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[4274] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[4275] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin2_
	HD[4276] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[4277] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[4278] = 32'b000111_01010_00000_0000000000001011; // beq 10 $zero _WhileExit2_
	HD[4279] = 32'b101101_00000000000000000000000100; // syscall 0
	HD[4280] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[4281] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[4282] = 32'b000001_11101_01100_0000000000000010; // lw 12 $fp 2
	HD[4283] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[4284] = 32'b000010_01011_01010_0000000000000000; // sw 10 11 0
	HD[4285] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[4286] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[4287] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[4288] = 32'b001011_00000000000000110001101000; // jump _WhileBegin2_
	HD[4289] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit2_
	HD[4290] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4291] = 32'b001111_11110_11111_0000000000000000; // push $ra / outputVector
	HD[4292] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[4293] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[4294] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin3_
	HD[4295] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[4296] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[4297] = 32'b000111_01010_00000_0000000000001011; // beq 10 $zero _WhileExit3_
	HD[4298] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[4299] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[4300] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[4301] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[4302] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[4303] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[4304] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[4305] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[4306] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[4307] = 32'b001011_00000000000000110001111011; // jump _WhileBegin3_
	HD[4308] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit3_
	HD[4309] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[4310] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0 / main
	HD[4311] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[4312] = 32'b000011_11101_11101_0000000000000001; // addi $fp $fp 1
	HD[4313] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[4314] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[4315] = 32'b001100_00000000000000110001100101; // jal inputVector
	HD[4316] = 32'b000100_11101_11101_0000000000000001; // subi $fp $fp 1
	HD[4317] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0
	HD[4318] = 32'b000101_00000_01011_0000000000000000; // li 11 0
	HD[4319] = 32'b000101_00000_01100_0000000000001010; // li 12 10
	HD[4320] = 32'b000011_11101_11101_0000000000000001; // addi $fp $fp 1
	HD[4321] = 32'b000010_11101_01100_0000000000000010; // sw 12 $fp 2
	HD[4322] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[4323] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[4324] = 32'b001100_00000000000000101111100001; // jal sort
	HD[4325] = 32'b000100_11101_11101_0000000000000001; // subi $fp $fp 1
	HD[4326] = 32'b101101_00000000000000000000000100; // syscall 0
	HD[4327] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[4328] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[4329] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0
	HD[4330] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[4331] = 32'b000001_11101_01100_0000000000000000; // lw 12 $fp 0
	HD[4332] = 32'b000011_11101_11101_0000000000000001; // addi $fp $fp 1
	HD[4333] = 32'b000010_11101_01100_0000000000000010; // sw 12 $fp 2
	HD[4334] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[4335] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[4336] = 32'b001100_00000000000000110001010011; // jal buscaBinaria
	HD[4337] = 32'b000100_11101_11101_0000000000000001; // subi $fp $fp 1
	HD[4338] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[4339] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[4340] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[4341] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0
	HD[4342] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[4343] = 32'b000011_11101_11101_0000000000000001; // addi $fp $fp 1
	HD[4344] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[4345] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[4346] = 32'b001100_00000000000000110001111000; // jal outputVector
	HD[4347] = 32'b000100_11101_11101_0000000000000001; // subi $fp $fp 1
	HD[4348] = 32'b101100_00000000000000000000001111; // return / _halt_

	/* Programa 03 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 5123> */
	HD[5123] = 32'b000011_11011_11101_0000000000001010; // addi $fp $global 10
	HD[5124] = 32'b001011_00000000000000101111101001; // jump main
	HD[5125] = 32'b001111_11110_11111_0000000000000000; // push $ra / mediaVector
	HD[5126] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[5127] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[5128] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[5129] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[5130] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin0_
	HD[5131] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[5132] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[5133] = 32'b000111_01010_00000_0000000000001100; // beq 10 $zero _WhileExit0_
	HD[5134] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3
	HD[5135] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[5136] = 32'b000001_11101_01100_0000000000000010; // lw 12 $fp 2
	HD[5137] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[5138] = 32'b000001_01011_01011_0000000000000000; // lw 11 11 0
	HD[5139] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[5140] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[5141] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[5142] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[5143] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[5144] = 32'b001011_00000000000000101110111111; // jump _WhileBegin0_
	HD[5145] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _WhileExit0_
	HD[5146] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[5147] = 32'b000000_01010_01011_01010_00000_001000; // div 10 10 11
	HD[5148] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[5149] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[5150] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[5151] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[5152] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[5153] = 32'b001111_11110_11111_0000000000000000; // push $ra / inputVector
	HD[5154] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[5155] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[5156] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin1_
	HD[5157] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[5158] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[5159] = 32'b000111_01010_00000_0000000000001011; // beq 10 $zero _WhileExit1_
	HD[5160] = 32'b101101_00000000000000000000000100; // syscall 0
	HD[5161] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[5162] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[5163] = 32'b000001_11101_01100_0000000000000010; // lw 12 $fp 2
	HD[5164] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[5165] = 32'b000010_01011_01010_0000000000000000; // sw 10 11 0
	HD[5166] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[5167] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[5168] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[5169] = 32'b001011_00000000000000101111011001; // jump _WhileBegin1_
	HD[5170] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit1_
	HD[5171] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[5172] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0 / main
	HD[5173] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[5174] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[5175] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[5176] = 32'b001100_00000000000000101111010110; // jal inputVector
	HD[5177] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0
	HD[5178] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[5179] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[5180] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[5181] = 32'b001100_00000000000000101110111010; // jal mediaVector
	HD[5182] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[5183] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[5184] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[5185] = 32'b101100_00000000000000000000001111; // return / _halt_

	/* Programa 04 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 6147> */
	HD[6147] = 32'b000011_11011_11101_0000000000001010; // addi $fp $global 10
	HD[6148] = 32'b001011_00000000000000110000010100; // jump main
	HD[6149] = 32'b001111_11110_11111_0000000000000000; // push $ra / mediaVector
	HD[6150] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[6151] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[6152] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[6153] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[6154] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin0_
	HD[6155] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[6156] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[6157] = 32'b000111_01010_00000_0000000000001100; // beq 10 $zero _WhileExit0_
	HD[6158] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3
	HD[6159] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[6160] = 32'b000001_11101_01100_0000000000000010; // lw 12 $fp 2
	HD[6161] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[6162] = 32'b000001_01011_01011_0000000000000000; // lw 11 11 0
	HD[6163] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[6164] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[6165] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[6166] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[6167] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[6168] = 32'b001011_00000000000000101110111111; // jump _WhileBegin0_
	HD[6169] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _WhileExit0_
	HD[6170] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[6171] = 32'b000000_01010_01011_01010_00000_001000; // div 10 10 11
	HD[6172] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[6173] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[6174] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[6175] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[6176] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[6177] = 32'b001111_11110_11111_0000000000000000; // push $ra / varianciaVector
	HD[6178] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[6179] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[6180] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[6181] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[6182] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[6183] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[6184] = 32'b000011_11101_11101_0000000000000110; // addi $fp $fp 6
	HD[6185] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[6186] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[6187] = 32'b001100_00000000000000101110111010; // jal mediaVector
	HD[6188] = 32'b000100_11101_11101_0000000000000110; // subi $fp $fp 6
	HD[6189] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[6190] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[6191] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin1_
	HD[6192] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[6193] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[6194] = 32'b000111_01010_00000_0000000000010010; // beq 10 $zero _WhileExit1_
	HD[6195] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[6196] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[6197] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[6198] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[6199] = 32'b000001_11101_01011_0000000000000100; // lw 11 $fp 4
	HD[6200] = 32'b000000_01010_01011_01010_00000_000110; // sub 10 10 11
	HD[6201] = 32'b000010_11101_01010_0000000000000101; // sw 10 $fp 5
	HD[6202] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3
	HD[6203] = 32'b000001_11101_01011_0000000000000101; // lw 11 $fp 5
	HD[6204] = 32'b000001_11101_01100_0000000000000101; // lw 12 $fp 5
	HD[6205] = 32'b000000_01011_01100_01011_00000_000111; // mult 11 11 12
	HD[6206] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[6207] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[6208] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[6209] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[6210] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[6211] = 32'b001011_00000000000000101111100100; // jump _WhileBegin1_
	HD[6212] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _WhileExit1_
	HD[6213] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[6214] = 32'b000000_01010_01011_01010_00000_001000; // div 10 10 11
	HD[6215] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[6216] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[6217] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[6218] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[6219] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[6220] = 32'b001111_11110_11111_0000000000000000; // push $ra / inputVector
	HD[6221] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[6222] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[6223] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin2_
	HD[6224] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[6225] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[6226] = 32'b000111_01010_00000_0000000000001011; // beq 10 $zero _WhileExit2_
	HD[6227] = 32'b101101_00000000000000000000000100; // syscall 0
	HD[6228] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[6229] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[6230] = 32'b000001_11101_01100_0000000000000010; // lw 12 $fp 2
	HD[6231] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[6232] = 32'b000010_01011_01010_0000000000000000; // sw 10 11 0
	HD[6233] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[6234] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[6235] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[6236] = 32'b001011_00000000000000110000000100; // jump _WhileBegin2_
	HD[6237] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit2_
	HD[6238] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[6239] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0 / main
	HD[6240] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[6241] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[6242] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[6243] = 32'b001100_00000000000000110000000001; // jal inputVector
	HD[6244] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0
	HD[6245] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[6246] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[6247] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[6248] = 32'b001100_00000000000000101111010110; // jal varianciaVector
	HD[6249] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[6250] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[6251] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[6252] = 32'b101100_00000000000000000000001111; // return / _halt_

	/* Programa 05 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 7171> */
	HD[7171] = 32'b000011_11011_11101_0000000000001010; // addi $fp $global 10
	HD[7172] = 32'b001011_00000000000000110000010000; // jump main
	HD[7173] = 32'b001111_11110_11111_0000000000000000; // push $ra / extremosVector
	HD[7174] = 32'b000101_00000_01010_0000000000000001; // li 10 1
	HD[7175] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[7176] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[7177] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[7178] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[7179] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[7180] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin0_
	HD[7181] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[7182] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[7183] = 32'b000111_01010_00000_0000000000011110; // beq 10 $zero _WhileExit0_
	HD[7184] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[7185] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[7186] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[7187] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[7188] = 32'b000001_11101_01011_0000000000000011; // lw 11 $fp 3
	HD[7189] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[7190] = 32'b000111_01010_00000_0000000000000111; // beq 10 $zero _ElseBegin0_
	HD[7191] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[7192] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[7193] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[7194] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[7195] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[7196] = 32'b001011_00000000000000101111011110; // jump _IfExit0_
	HD[7197] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0 / _ElseBegin0_
	HD[7198] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[7199] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[7200] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[7201] = 32'b000001_11101_01011_0000000000000100; // lw 11 $fp 4
	HD[7202] = 32'b000000_01010_01011_01010_00000_010010; // sgt 10 10 11
	HD[7203] = 32'b000111_01010_00000_0000000000000110; // beq 10 $zero _IfExit1_
	HD[7204] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[7205] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[7206] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[7207] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[7208] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[7209] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _IfExit1_ _IfExit0_
	HD[7210] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[7211] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[7212] = 32'b001011_00000000000000101111000001; // jump _WhileBegin0_
	HD[7213] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _WhileExit0_
	HD[7214] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[7215] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[7216] = 32'b000001_11101_01010_0000000000000100; // lw 10 $fp 4
	HD[7217] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[7218] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[7219] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[7220] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[7221] = 32'b001111_11110_11111_0000000000000000; // push $ra / inputVector
	HD[7222] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[7223] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[7224] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin1_
	HD[7225] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[7226] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[7227] = 32'b000111_01010_00000_0000000000001011; // beq 10 $zero _WhileExit1_
	HD[7228] = 32'b101101_00000000000000000000000100; // syscall 0
	HD[7229] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[7230] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[7231] = 32'b000001_11101_01100_0000000000000010; // lw 12 $fp 2
	HD[7232] = 32'b000000_01011_01100_01011_00000_000101; // add 11 11 12
	HD[7233] = 32'b000010_01011_01010_0000000000000000; // sw 10 11 0
	HD[7234] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[7235] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[7236] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[7237] = 32'b001011_00000000000000101111101101; // jump _WhileBegin1_
	HD[7238] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit1_
	HD[7239] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[7240] = 32'b001111_11110_11111_0000000000000000; // push $ra / outputVector
	HD[7241] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[7242] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[7243] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin2_
	HD[7244] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[7245] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[7246] = 32'b000111_01010_00000_0000000000001011; // beq 10 $zero _WhileExit2_
	HD[7247] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[7248] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[7249] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[7250] = 32'b000001_01010_01010_0000000000000000; // lw 10 10 0
	HD[7251] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[7252] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[7253] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[7254] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[7255] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[7256] = 32'b001011_00000000000000110000000000; // jump _WhileBegin2_
	HD[7257] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit2_
	HD[7258] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[7259] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0 / main
	HD[7260] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[7261] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[7262] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[7263] = 32'b001100_00000000000000101111101010; // jal inputVector
	HD[7264] = 32'b000011_11011_01010_0000000000000000; // addi 10 $global 0
	HD[7265] = 32'b000101_00000_01011_0000000000001010; // li 11 10
	HD[7266] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[7267] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[7268] = 32'b001100_00000000000000101110111010; // jal extremosVector
	HD[7269] = 32'b101100_00000000000000000000001111; // return / _halt_

	/* Programa 06 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 8195> */
	HD[8195] = 32'b000011_11011_11101_0000000000000000; // addi $fp $global 0
	HD[8196] = 32'b001011_00000000000000101111010111; // jump main
	HD[8197] = 32'b001111_11110_11111_0000000000000000; // push $ra / gcd
	HD[8198] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1
	HD[8199] = 32'b000101_00000_01011_0000000000000000; // li 11 0
	HD[8200] = 32'b000000_01010_01011_01010_00000_010011; // set 10 10 11
	HD[8201] = 32'b000111_01010_00000_0000000000000110; // beq 10 $zero _ElseBegin0_
	HD[8202] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[8203] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[8204] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[8205] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[8206] = 32'b001011_00000000000000101111010101; // jump _IfExit0_
	HD[8207] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1 / _ElseBegin0_
	HD[8208] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[8209] = 32'b000001_11101_01100_0000000000000000; // lw 12 $fp 0
	HD[8210] = 32'b000001_11101_01101_0000000000000001; // lw 13 $fp 1
	HD[8211] = 32'b000000_01100_01101_01100_00000_001000; // div 12 12 13
	HD[8212] = 32'b000001_11101_01101_0000000000000001; // lw 13 $fp 1
	HD[8213] = 32'b000000_01100_01101_01100_00000_000111; // mult 12 12 13
	HD[8214] = 32'b000000_01011_01100_01011_00000_000110; // sub 11 11 12
	HD[8215] = 32'b000011_11101_11101_0000000000000010; // addi $fp $fp 2
	HD[8216] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[8217] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[8218] = 32'b001100_00000000000000101110111010; // jal gcd
	HD[8219] = 32'b000100_11101_11101_0000000000000010; // subi $fp $fp 2
	HD[8220] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[8221] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[8222] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[8223] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[8224] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit0_
	HD[8225] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[8226] = 32'b101101_00000000000000000000000100; // syscall 0 / main
	HD[8227] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[8228] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[8229] = 32'b101101_00000000000000000000000100; // syscall 0
	HD[8230] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[8231] = 32'b000010_11101_01010_0000000000000001; // sw 10 $fp 1
	HD[8232] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[8233] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[8234] = 32'b000011_11101_11101_0000000000000010; // addi $fp $fp 2
	HD[8235] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[8236] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[8237] = 32'b001100_00000000000000101110111010; // jal gcd
	HD[8238] = 32'b000100_11101_11101_0000000000000010; // subi $fp $fp 2
	HD[8239] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[8240] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[8241] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[8242] = 32'b101100_00000000000000000000001111; // return / _halt_

	/* Programa 07 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 9219> */
	HD[9219] = 32'b000011_11011_11101_0000000000000000; // addi $fp $global 0
	HD[9220] = 32'b001011_00000000000000101111100111; // jump main
	HD[9221] = 32'b001111_11110_11111_0000000000000000; // push $ra / fibonacci
	HD[9222] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[9223] = 32'b000101_00000_01011_0000000000000000; // li 11 0
	HD[9224] = 32'b000000_01010_01011_01010_00000_010010; // sgt 10 10 11
	HD[9225] = 32'b000000_01010_00000_01010_00000_010011; // set 10 10 $zero
	HD[9226] = 32'b000111_01010_00000_0000000000000101; // beq 10 $zero _ElseBegin0_
	HD[9227] = 32'b000101_00000_11100_0000000000000000; // li $rv 0
	HD[9228] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[9229] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[9230] = 32'b001011_00000000000000101111100101; // jump _IfExit0_
	HD[9231] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0 / _ElseBegin0_
	HD[9232] = 32'b000101_00000_01011_0000000000000001; // li 11 1
	HD[9233] = 32'b000000_01010_01011_01010_00000_010011; // set 10 10 11
	HD[9234] = 32'b000111_01010_00000_0000000000000101; // beq 10 $zero _ElseBegin1_
	HD[9235] = 32'b000101_00000_11100_0000000000000001; // li $rv 1
	HD[9236] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[9237] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[9238] = 32'b001011_00000000000000101111100101; // jump _IfExit1_
	HD[9239] = 32'b000101_00000_01010_0000000000000000; // li 10 0 / _ElseBegin1_
	HD[9240] = 32'b000010_11101_01010_0000000000000001; // sw 10 $fp 1
	HD[9241] = 32'b000101_00000_01010_0000000000000001; // li 10 1
	HD[9242] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[9243] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[9244] = 32'b000001_11101_01010_0000000000000100; // lw 10 $fp 4 / _WhileBegin0_
	HD[9245] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[9246] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[9247] = 32'b000111_01010_00000_0000000000001101; // beq 10 $zero _WhileExit0_
	HD[9248] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[9249] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[9250] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[9251] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[9252] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[9253] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[9254] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3
	HD[9255] = 32'b000010_11101_01010_0000000000000001; // sw 10 $fp 1
	HD[9256] = 32'b000001_11101_01010_0000000000000100; // lw 10 $fp 4
	HD[9257] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[9258] = 32'b000010_11101_01010_0000000000000100; // sw 10 $fp 4
	HD[9259] = 32'b001011_00000000000000101111010001; // jump _WhileBegin0_
	HD[9260] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileExit0_
	HD[9261] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[9262] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[9263] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[9264] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit1_ _IfExit0_
	HD[9265] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[9266] = 32'b101101_00000000000000000000000100; // syscall 0 / main
	HD[9267] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[9268] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[9269] = 32'b001100_00000000000000101110111010; // jal fibonacci
	HD[9270] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[9271] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[9272] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[9273] = 32'b101100_00000000000000000000001111; // return / _halt_

	/* Programa 08 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 10243> */
	HD[10243] = 32'b000011_11011_11101_0000000000000000; // addi $fp $global 0
	HD[10244] = 32'b001011_00000000000000101111010001; // jump main
	HD[10245] = 32'b001111_11110_11111_0000000000000000; // push $ra / fatorial
	HD[10246] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[10247] = 32'b000101_00000_01011_0000000000000010; // li 11 2
	HD[10248] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[10249] = 32'b000111_01010_00000_0000000000000101; // beq 10 $zero _ElseBegin0_
	HD[10250] = 32'b000101_00000_11100_0000000000000001; // li $rv 1
	HD[10251] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[10252] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[10253] = 32'b001011_00000000000000101111001111; // jump _IfExit0_
	HD[10254] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0 / _ElseBegin0_
	HD[10255] = 32'b000100_01010_01010_0000000000000001; // subi 10 10 1
	HD[10256] = 32'b000011_11101_11101_0000000000000001; // addi $fp $fp 1
	HD[10257] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[10258] = 32'b001100_00000000000000101110111010; // jal fatorial
	HD[10259] = 32'b000100_11101_11101_0000000000000001; // subi $fp $fp 1
	HD[10260] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[10261] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[10262] = 32'b000000_01010_01011_01010_00000_000111; // mult 10 10 11
	HD[10263] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[10264] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[10265] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[10266] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit0_
	HD[10267] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[10268] = 32'b101101_00000000000000000000000100; // syscall 0 / main
	HD[10269] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[10270] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[10271] = 32'b001100_00000000000000101110111010; // jal fatorial
	HD[10272] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[10273] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[10274] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[10275] = 32'b101100_00000000000000000000001111; // return / _halt_

	/* Programa 09 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 11267> */
	HD[11267] = 32'b000011_11011_11101_0000000000000000; // addi $fp $global 0
	HD[11268] = 32'b001011_00000000000000110000001000; // jump main
	HD[11269] = 32'b001111_11110_11111_0000000000000000; // push $ra / calculadora
	HD[11270] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[11271] = 32'b000101_00000_01011_0000000000000001; // li 11 1
	HD[11272] = 32'b000000_01010_01011_01010_00000_010011; // set 10 10 11
	HD[11273] = 32'b000111_01010_00000_0000000000001000; // beq 10 $zero _ElseBegin0_
	HD[11274] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[11275] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[11276] = 32'b000000_01010_01011_01010_00000_000101; // add 10 10 11
	HD[11277] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[11278] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[11279] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[11280] = 32'b001011_00000000000000110000000110; // jump _IfExit0_
	HD[11281] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _ElseBegin0_
	HD[11282] = 32'b000101_00000_01011_0000000000000010; // li 11 2
	HD[11283] = 32'b000000_01010_01011_01010_00000_010011; // set 10 10 11
	HD[11284] = 32'b000111_01010_00000_0000000000001000; // beq 10 $zero _ElseBegin1_
	HD[11285] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[11286] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[11287] = 32'b000000_01010_01011_01010_00000_000110; // sub 10 10 11
	HD[11288] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[11289] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[11290] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[11291] = 32'b001011_00000000000000110000000110; // jump _IfExit1_
	HD[11292] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _ElseBegin1_
	HD[11293] = 32'b000101_00000_01011_0000000000000011; // li 11 3
	HD[11294] = 32'b000000_01010_01011_01010_00000_010011; // set 10 10 11
	HD[11295] = 32'b000111_01010_00000_0000000000001000; // beq 10 $zero _ElseBegin2_
	HD[11296] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[11297] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[11298] = 32'b000000_01010_01011_01010_00000_000111; // mult 10 10 11
	HD[11299] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[11300] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[11301] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[11302] = 32'b001011_00000000000000110000000110; // jump _IfExit2_
	HD[11303] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _ElseBegin2_
	HD[11304] = 32'b000101_00000_01011_0000000000000100; // li 11 4
	HD[11305] = 32'b000000_01010_01011_01010_00000_010011; // set 10 10 11
	HD[11306] = 32'b000111_01010_00000_0000000000001000; // beq 10 $zero _ElseBegin3_
	HD[11307] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[11308] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[11309] = 32'b000000_01010_01011_01010_00000_001000; // div 10 10 11
	HD[11310] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[11311] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[11312] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[11313] = 32'b001011_00000000000000110000000110; // jump _IfExit3_
	HD[11314] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _ElseBegin3_
	HD[11315] = 32'b000101_00000_01011_0000000000000101; // li 11 5
	HD[11316] = 32'b000000_01010_01011_01010_00000_010011; // set 10 10 11
	HD[11317] = 32'b000111_01010_00000_0000000000001100; // beq 10 $zero _ElseBegin4_
	HD[11318] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[11319] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[11320] = 32'b000001_11101_01100_0000000000000001; // lw 12 $fp 1
	HD[11321] = 32'b000000_01011_01100_01011_00000_001000; // div 11 11 12
	HD[11322] = 32'b000001_11101_01100_0000000000000001; // lw 12 $fp 1
	HD[11323] = 32'b000000_01011_01100_01011_00000_000111; // mult 11 11 12
	HD[11324] = 32'b000000_01010_01011_01010_00000_000110; // sub 10 10 11
	HD[11325] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[11326] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[11327] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[11328] = 32'b001011_00000000000000110000000110; // jump _IfExit4_
	HD[11329] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _ElseBegin4_
	HD[11330] = 32'b000101_00000_01011_0000000000000110; // li 11 6
	HD[11331] = 32'b000000_01010_01011_01010_00000_010011; // set 10 10 11
	HD[11332] = 32'b000111_01010_00000_0000000000001010; // beq 10 $zero _ElseBegin5_
	HD[11333] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[11334] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[11335] = 32'b000000_01010_01011_01010_00000_000111; // mult 10 10 11
	HD[11336] = 32'b000101_00000_01011_0000000001100100; // li 11 100
	HD[11337] = 32'b000000_01010_01011_01010_00000_001000; // div 10 10 11
	HD[11338] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[11339] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[11340] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[11341] = 32'b001011_00000000000000110000000110; // jump _IfExit5_
	HD[11342] = 32'b000101_00000_11100_0000000000000000; // li $rv 0 / _ElseBegin5_
	HD[11343] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[11344] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[11345] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit5_ _IfExit4_ _IfExit3_ _IfExit2_ _IfExit1_ _IfExit0_
	HD[11346] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[11347] = 32'b101101_00000000000000000000000100; // syscall 0 / main
	HD[11348] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[11349] = 32'b000010_11101_01010_0000000000000001; // sw 10 $fp 1
	HD[11350] = 32'b101101_00000000000000000000000100; // syscall 0
	HD[11351] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[11352] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[11353] = 32'b101101_00000000000000000000000100; // syscall 0
	HD[11354] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[11355] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[11356] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1
	HD[11357] = 32'b000001_11101_01011_0000000000000010; // lw 11 $fp 2
	HD[11358] = 32'b000001_11101_01100_0000000000000011; // lw 12 $fp 3
	HD[11359] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
	HD[11360] = 32'b000010_11101_01100_0000000000000010; // sw 12 $fp 2
	HD[11361] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[11362] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[11363] = 32'b001100_00000000000000101110111010; // jal calculadora
	HD[11364] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
	HD[11365] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[11366] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[11367] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[11368] = 32'b101100_00000000000000000000001111; // return / _halt_

	/* Programa 10 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 12291> */
	HD[12291] = 32'b000011_11011_11101_0000000000000000; // addi $fp $global 0
	HD[12292] = 32'b001011_00000000000000101111101001; // jump main
	HD[12293] = 32'b001111_11110_11111_0000000000000000; // push $ra / potencia
	HD[12294] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1
	HD[12295] = 32'b000101_00000_01011_0000000000000000; // li 11 0
	HD[12296] = 32'b000000_01010_01011_01010_00000_010011; // set 10 10 11
	HD[12297] = 32'b000111_01010_00000_0000000000000101; // beq 10 $zero _ElseBegin0_
	HD[12298] = 32'b000101_00000_11100_0000000000000001; // li $rv 1
	HD[12299] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[12300] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[12301] = 32'b001011_00000000000000101111100111; // jump _IfExit0_
	HD[12302] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0 / _ElseBegin0_
	HD[12303] = 32'b000101_00000_01011_0000000000000000; // li 11 0
	HD[12304] = 32'b000000_01010_01011_01010_00000_010011; // set 10 10 11
	HD[12305] = 32'b000111_01010_00000_0000000000000101; // beq 10 $zero _ElseBegin1_
	HD[12306] = 32'b000101_00000_11100_0000000000000000; // li $rv 0
	HD[12307] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[12308] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[12309] = 32'b001011_00000000000000101111100111; // jump _IfExit1_
	HD[12310] = 32'b000001_11101_01010_0000000000000001; // lw 10 $fp 1 / _ElseBegin1_
	HD[12311] = 32'b000101_00000_01011_0000000000000000; // li 11 0
	HD[12312] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[12313] = 32'b000111_01010_00000_0000000000000101; // beq 10 $zero _ElseBegin2_
	HD[12314] = 32'b000101_00000_11100_0000000000000000; // li $rv 0
	HD[12315] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[12316] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[12317] = 32'b001011_00000000000000101111100111; // jump _IfExit2_
	HD[12318] = 32'b000101_00000_01010_0000000000000001; // li 10 1 / _ElseBegin2_
	HD[12319] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[12320] = 32'b000101_00000_01010_0000000000000000; // li 10 0
	HD[12321] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[12322] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2 / _WhileBegin0_
	HD[12323] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[12324] = 32'b000000_01010_01011_01010_00000_010001; // slt 10 10 11
	HD[12325] = 32'b000111_01010_00000_0000000000001001; // beq 10 $zero _WhileExit0_
	HD[12326] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3
	HD[12327] = 32'b000001_11101_01011_0000000000000000; // lw 11 $fp 0
	HD[12328] = 32'b000000_01010_01011_01010_00000_000111; // mult 10 10 11
	HD[12329] = 32'b000010_11101_01010_0000000000000011; // sw 10 $fp 3
	HD[12330] = 32'b000001_11101_01010_0000000000000010; // lw 10 $fp 2
	HD[12331] = 32'b000011_01010_01010_0000000000000001; // addi 10 10 1
	HD[12332] = 32'b000010_11101_01010_0000000000000010; // sw 10 $fp 2
	HD[12333] = 32'b001011_00000000000000101111010111; // jump _WhileBegin0_
	HD[12334] = 32'b000001_11101_01010_0000000000000011; // lw 10 $fp 3 / _WhileExit0_
	HD[12335] = 32'b000000_01010_11100_00000_00000_010000; // move $rv 10
	HD[12336] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[12337] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[12338] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit2_ _IfExit1_ _IfExit0_
	HD[12339] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[12340] = 32'b101101_00000000000000000000000100; // syscall 0 / main
	HD[12341] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[12342] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[12343] = 32'b101101_00000000000000000000000100; // syscall 0
	HD[12344] = 32'b000000_11001_01010_00000_00000_010000; // move 10 25
	HD[12345] = 32'b000010_11101_01010_0000000000000001; // sw 10 $fp 1
	HD[12346] = 32'b000001_11101_01010_0000000000000000; // lw 10 $fp 0
	HD[12347] = 32'b000001_11101_01011_0000000000000001; // lw 11 $fp 1
	HD[12348] = 32'b000011_11101_11101_0000000000000010; // addi $fp $fp 2
	HD[12349] = 32'b000010_11101_01011_0000000000000001; // sw 11 $fp 1
	HD[12350] = 32'b000010_11101_01010_0000000000000000; // sw 10 $fp 0
	HD[12351] = 32'b001100_00000000000000101110111010; // jal potencia
	HD[12352] = 32'b000100_11101_11101_0000000000000010; // subi $fp $fp 2
	HD[12353] = 32'b000000_11100_01010_00000_00000_010000; // move 10 $rv
	HD[12354] = 32'b000000_01010_11001_00000_00000_010000; // move 25 10
	HD[12355] = 32'b101101_00000000000000000000001000; // syscall 1
	HD[12356] = 32'b101100_00000000000000000000001111; // return / _halt_
	
	/* Programa 11 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 13315> */
	HD[13315] = 32'b000101_00000_00001_0000000000000111; // li 1 7
	HD[13316] = 32'b010001_00001_00000_0000000000000000; // send 1
	HD[13317] = 32'b000101_00000_00010_0000000000001010; // li 2 10
	HD[13318] = 32'b000101_00000_00100_0000000000001100; // li 4 12
	HD[13319] = 32'b001010_00001_00000_0000000000000000; // out 1
	HD[13320] = 32'b010010_00000_00101_0000000000000000; // recv 5
	HD[13321] = 32'b001010_00101_00000_0000000000000000; // out 5
	HD[13322] = 32'b101100_00000000000000000000001111; // return
	
	/* Programa 12 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 14339> */
	HD[14339] = 32'b000101_00000_00001_0000000000000111; // li 1 7
	HD[14340] = 32'b001010_00001_00000_0000000000000000; // out 1
	HD[14341] = 32'b010010_00000_00101_0000000000000000; // recv 5
	HD[14342] = 32'b001010_00101_00000_0000000000000000; // out 5
	HD[14343] = 32'b000011_00101_00101_0000000000001010; // addi 5 10
	HD[14344] = 32'b010001_00101_00000_0000000000000000; // send 5
	HD[14345] = 32'b001010_00101_00000_0000000000000000; // out 5
	HD[14346] = 32'b101100_00000000000000000000001111; // return
	
	/* Programa 13 */
	/* Parameters: <mem_offset = 3000> <priority_system = false> <index_begin = 15363> */
	HD[15363] = 32'b000101_00000_11011_0000000000000000; // li $global 0
	HD[15364] = 32'b000011_11011_11101_0000000000000000; // addi $fp $global 0
	HD[15365] = 32'b001011_00000000000000110000100111; // jump main
	HD[15366] = 32'b001111_11110_11111_0000000000000000; // push $ra / sleep
	HD[15367] = 32'b000101_00000_00010_0000000000000000; // li 2 0
	HD[15368] = 32'b000010_11101_00010_0000000000000001; // sw 2 $fp 1
	HD[15369] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
	HD[15370] = 32'b000101_00000_00011_0000000000011001; // li 3 25
	HD[15371] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[15372] = 32'b000101_00000_00011_0000000000000100; // li 3 4
	HD[15373] = 32'b000000_00010_00011_00010_00000_001000; // div 2 2 3
	HD[15374] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
	HD[15375] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1 / _WhileBegin0_
	HD[15376] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
	HD[15377] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[15378] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _WhileExit0_
	HD[15379] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1
	HD[15380] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
	HD[15381] = 32'b000010_11101_00010_0000000000000001; // sw 2 $fp 1
	HD[15382] = 32'b001011_00000000000000101111000100; // jump _WhileBegin0_
	HD[15383] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit0_
	HD[15384] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[15385] = 32'b001111_11110_11111_0000000000000000; // push $ra / mod
	HD[15386] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
	HD[15387] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
	HD[15388] = 32'b000001_11101_00100_0000000000000001; // lw 4 $fp 1
	HD[15389] = 32'b000000_00011_00100_00011_00000_001000; // div 3 3 4
	HD[15390] = 32'b000001_11101_00100_0000000000000001; // lw 4 $fp 1
	HD[15391] = 32'b000000_00011_00100_00011_00000_000111; // mult 3 3 4
	HD[15392] = 32'b000000_00010_00011_00010_00000_000110; // sub 2 2 3
	HD[15393] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
	HD[15394] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[15395] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[15396] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[15397] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[15398] = 32'b001111_11110_11111_0000000000000000; // push $ra / print_value
	HD[15399] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
	HD[15400] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[15401] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
	HD[15402] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
	HD[15403] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
	HD[15404] = 32'b001100_00000000000000101111001110; // jal mod
	HD[15405] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
	HD[15406] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
	HD[15407] = 32'b000011_00010_00010_0000000000110000; // addi 2 2 48
	HD[15408] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
	HD[15409] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1
	HD[15410] = 32'b000101_00000_00011_0000000000010000; // li 3 16
	HD[15411] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[15412] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
	HD[15413] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[15414] = 32'b000001_11101_00011_0000000000000011; // lw 3 $fp 3
	HD[15415] = 32'b100111_00010_00011_00011_00000000000; // lcdwrite 2 3 3
	HD[15416] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
	HD[15417] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[15418] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[15419] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[15420] = 32'b000111_00010_00000_0000000000001110; // beq 2 $zero _ElseBegin0_
	HD[15421] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
	HD[15422] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[15423] = 32'b000000_00010_00011_00010_00000_001000; // div 2 2 3
	HD[15424] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[15425] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
	HD[15426] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
	HD[15427] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
	HD[15428] = 32'b001100_00000000000000101111001110; // jal mod
	HD[15429] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
	HD[15430] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
	HD[15431] = 32'b000011_00010_00010_0000000000110000; // addi 2 2 48
	HD[15432] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
	HD[15433] = 32'b001011_00000000000000110000000001; // jump _IfExit0_
	HD[15434] = 32'b000101_00000_00010_0000000000100000; // li 2 32 / _ElseBegin0_
	HD[15435] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
	HD[15436] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1 / _IfExit0_
	HD[15437] = 32'b000101_00000_00011_0000000000010000; // li 3 16
	HD[15438] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[15439] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
	HD[15440] = 32'b000100_00011_00011_0000000000000001; // subi 3 3 1
	HD[15441] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[15442] = 32'b000001_11101_00011_0000000000000011; // lw 3 $fp 3
	HD[15443] = 32'b100111_00010_00011_00011_00000000000; // lcdwrite 2 3 3
	HD[15444] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
	HD[15445] = 32'b000101_00000_00011_0000000001100100; // li 3 100
	HD[15446] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
	HD[15447] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
	HD[15448] = 32'b000111_00010_00000_0000000000001110; // beq 2 $zero _ElseBegin1_
	HD[15449] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
	HD[15450] = 32'b000101_00000_00011_0000000001100100; // li 3 100
	HD[15451] = 32'b000000_00010_00011_00010_00000_001000; // div 2 2 3
	HD[15452] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[15453] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
	HD[15454] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
	HD[15455] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
	HD[15456] = 32'b001100_00000000000000101111001110; // jal mod
	HD[15457] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
	HD[15458] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
	HD[15459] = 32'b000011_00010_00010_0000000000110000; // addi 2 2 48
	HD[15460] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
	HD[15461] = 32'b001011_00000000000000110000011101; // jump _IfExit1_
	HD[15462] = 32'b000101_00000_00010_0000000000100000; // li 2 32 / _ElseBegin1_
	HD[15463] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
	HD[15464] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1 / _IfExit1_
	HD[15465] = 32'b000101_00000_00011_0000000000010000; // li 3 16
	HD[15466] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
	HD[15467] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
	HD[15468] = 32'b000100_00011_00011_0000000000000010; // subi 3 3 2
	HD[15469] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
	HD[15470] = 32'b000001_11101_00011_0000000000000011; // lw 3 $fp 3
	HD[15471] = 32'b100111_00010_00011_00011_00000000000; // lcdwrite 2 3 3
	HD[15472] = 32'b010000_11110_11111_0000000000000000; // pop $ra
	HD[15473] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
	HD[15474] = 32'b100110_00000000000000000000000000; // lcdclean / main
	HD[15475] = 32'b100111_00001_00000_00000_00001010110; // lcdwrite 1 86
	HD[15476] = 32'b100111_00010_00000_00000_00001100001; // lcdwrite 2 97
	HD[15477] = 32'b100111_00011_00000_00000_00001101100; // lcdwrite 3 108
	HD[15478] = 32'b100111_00100_00000_00000_00001101111; // lcdwrite 4 111
	HD[15479] = 32'b100111_00101_00000_00000_00001110010; // lcdwrite 5 114
	HD[15480] = 32'b100111_00110_00000_00000_00000111010; // lcdwrite 6 58
	HD[15481] = 32'b100111_10001_00000_00000_00001000110; // lcdwrite 17 70
	HD[15482] = 32'b100111_10010_00000_00000_00001010000; // lcdwrite 18 80
	HD[15483] = 32'b100111_10011_00000_00000_00001000111; // lcdwrite 19 71
	HD[15484] = 32'b100111_10100_00000_00000_00001000001; // lcdwrite 20 65
	HD[15485] = 32'b100111_10110_00000_00000_00001010011; // lcdwrite 22 83
	HD[15486] = 32'b100111_10111_00000_00000_00001001111; // lcdwrite 23 79
	HD[15487] = 32'b100111_11001_00000_00000_00001010011; // lcdwrite 25 83
	HD[15488] = 32'b100111_11010_00000_00000_00001001100; // lcdwrite 26 76
	HD[15489] = 32'b100111_11011_00000_00000_00001000001; // lcdwrite 27 65
	HD[15490] = 32'b100111_11100_00000_00000_00001010110; // lcdwrite 28 86
	HD[15491] = 32'b100111_11101_00000_00000_00001000101; // lcdwrite 29 69
	HD[15492] = 32'b000101_00000_00010_0000000000000001; // li 2 1 / _WhileBegin1_
	HD[15493] = 32'b000111_00010_00000_0000000000011100; // beq 2 $zero _WhileExit1_
	HD[15494] = 32'b010010_00000_00010_0000000000000000; // recv 2
	HD[15495] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
	HD[15496] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
	HD[15497] = 32'b000101_00000_00011_0000000000001010; // li 3 10
	HD[15498] = 32'b000011_11101_11101_0000000000000001; // addi $fp $fp 1
	HD[15499] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
	HD[15500] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
	HD[15501] = 32'b001100_00000000000000101111001110; // jal mod
	HD[15502] = 32'b000100_11101_11101_0000000000000001; // subi $fp $fp 1
	HD[15503] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
	HD[15504] = 32'b100111_01110_00010_00010_00000000000; // lcdwrite 14 2 2
	HD[15505] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
	HD[15506] = 32'b000101_00000_00011_0000000000000000; // li 3 0
	HD[15507] = 32'b000101_00000_00100_0000000000001101; // li 4 13
	HD[15508] = 32'b000011_11101_11101_0000000000000001; // addi $fp $fp 1
	HD[15509] = 32'b000010_11101_00100_0000000000000010; // sw 4 $fp 2
	HD[15510] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
	HD[15511] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
	HD[15512] = 32'b001100_00000000000000101111011011; // jal print_value
	HD[15513] = 32'b000100_11101_11101_0000000000000001; // subi $fp $fp 1
	HD[15514] = 32'b100111_01101_00000_00000_00000101100; // lcdwrite 13 44
	HD[15515] = 32'b000101_00000_00010_0000000001100100; // li 2 100
	HD[15516] = 32'b000011_11101_11101_0000000000000001; // addi $fp $fp 1
	HD[15517] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
	HD[15518] = 32'b001100_00000000000000101110111011; // jal sleep
	HD[15519] = 32'b000100_11101_11101_0000000000000001; // subi $fp $fp 1
	HD[15520] = 32'b001011_00000000000000110000111001; // jump _WhileBegin1_
	HD[15521] = 32'b100110_00000000000000000000000000; // lcdclean / _WhileExit1_
	HD[15522] = 32'b11111111111111111111111111111111; // halt / _halt_
	end 
	
	always @ (posedge write_clock)
	begin
		if (hdWrite == 1'b1) begin
			HD[trilha*HD_SETORES_SIZE+setor] <= data;
		end
	end
	
	always @ (posedge read_clock)
	begin
		dataRead <= HD[trilha*HD_SETORES_SIZE+setor];
	end
	
	assign dataOut = (hdRead == 1'b1) ? dataRead : 0;
	
	/*initial begin
		HD[0][0] <= 32'b000101_00000_00010_0000000011001000; // li 2 200
		HD[0][1] <= 32'b001010_00010_00000_0000000000000000; // out 2
		HD[0][2] <= 32'b11111111111111111111111111111111; // halt
	end*/
	
endmodule 
module ram_inst(write_clock, read_clock, reset, instWrite, addr, datain, memAddress, out);
	
	parameter DATA_WIDTH = 32; // X bits 
	parameter RAM_BITS = 12; // X instructions
	localparam RAM_SIZE = 2**RAM_BITS; 
	
	input write_clock, read_clock, reset, instWrite;
	input [DATA_WIDTH-1:0] addr, memAddress;  
	input [DATA_WIDTH-1:0] datain;
	output reg [DATA_WIDTH-1:0] out;
	
	reg [DATA_WIDTH-1:0] RAM_INST [RAM_SIZE-1:0]; // RAM_SIZE words of 32-bit memory
	
	initial 
	begin : INIT
	
		
		//RAM_INST[2] = 32'b000101_00000_00010_0000000000000101; // li 2 5
		//RAM_INST[3] = 32'b100101_00000_00010_00001_00000_000000; // regtohd 0 2 1
		//RAM_INST[4] = 32'b100100_00000_00010_00011_00000_000000; // hdtoreg 0 2 3
		//RAM_INST[5] = 32'b001010_00011_00000_0000000000000000; // out 3
        //RAM_INST[0] = 32'b001010_00000_00000_0000000000000000; // out 0
        //RAM_INST[1] = 32'b111111_00000_00000_0000000000000000; // halt
	end 
	
	always @ (posedge write_clock)
	begin
	
		if (instWrite) begin 
			RAM_INST[addr] <= datain;
		end
		
		if (reset) begin
		/*
			RAM_INST[0] = 32'b000101_00000_11011_0000000000000000; // li $global 0
RAM_INST[1] = 32'b000011_11011_11101_0000000000001010; // addi $fp $global 10
RAM_INST[2] = 32'b001011_00000000000000000111001011; // jump main
RAM_INST[3] = 32'b001111_11110_11111_0000000000000000; // push $ra / minloc
RAM_INST[4] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1
RAM_INST[5] = 32'b000010_11101_00010_0000000000000101; // sw 2 $fp 5
RAM_INST[6] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[7] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[8] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[9] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[10] = 32'b000010_11101_00010_0000000000000100; // sw 2 $fp 4
RAM_INST[11] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1
RAM_INST[12] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
RAM_INST[13] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
RAM_INST[14] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3 / _WhileBegin0_
RAM_INST[15] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
RAM_INST[16] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[17] = 32'b000111_00010_00000_0000000000010011; // beq 2 $zero _WhileExit0_
RAM_INST[18] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[19] = 32'b000001_11101_00011_0000000000000011; // lw 3 $fp 3
RAM_INST[20] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[21] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[22] = 32'b000001_11101_00011_0000000000000100; // lw 3 $fp 4
RAM_INST[23] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[24] = 32'b000111_00010_00000_0000000000001000; // beq 2 $zero _IfExit0_
RAM_INST[25] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[26] = 32'b000001_11101_00011_0000000000000011; // lw 3 $fp 3
RAM_INST[27] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[28] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[29] = 32'b000010_11101_00010_0000000000000100; // sw 2 $fp 4
RAM_INST[30] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3
RAM_INST[31] = 32'b000010_11101_00010_0000000000000101; // sw 2 $fp 5
RAM_INST[32] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3 / _IfExit0_
RAM_INST[33] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
RAM_INST[34] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
RAM_INST[35] = 32'b001011_00000000000000000000001110; // jump _WhileBegin0_
RAM_INST[36] = 32'b000001_11101_00010_0000000000000101; // lw 2 $fp 5 / _WhileExit0_
RAM_INST[37] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[38] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[39] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[40] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[41] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[42] = 32'b001111_11110_11111_0000000000000000; // push $ra / sort
RAM_INST[43] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1
RAM_INST[44] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
RAM_INST[45] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3 / _WhileBegin1_
RAM_INST[46] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
RAM_INST[47] = 32'b000100_00011_00011_0000000000000001; // subi 3 3 1
RAM_INST[48] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[49] = 32'b000111_00010_00000_0000000000100010; // beq 2 $zero _WhileExit1_
RAM_INST[50] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[51] = 32'b000001_11101_00011_0000000000000011; // lw 3 $fp 3
RAM_INST[52] = 32'b000001_11101_00100_0000000000000010; // lw 4 $fp 2
RAM_INST[53] = 32'b000011_11101_11101_0000000000000110; // addi $fp $fp 6
RAM_INST[54] = 32'b000010_11101_00100_0000000000000010; // sw 4 $fp 2
RAM_INST[55] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[56] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[57] = 32'b001100_00000000000000000000000011; // jal minloc
RAM_INST[58] = 32'b000100_11101_11101_0000000000000110; // subi $fp $fp 6
RAM_INST[59] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[60] = 32'b000010_11101_00010_0000000000000100; // sw 2 $fp 4
RAM_INST[61] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[62] = 32'b000001_11101_00011_0000000000000100; // lw 3 $fp 4
RAM_INST[63] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[64] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[65] = 32'b000010_11101_00010_0000000000000101; // sw 2 $fp 5
RAM_INST[66] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[67] = 32'b000001_11101_00011_0000000000000011; // lw 3 $fp 3
RAM_INST[68] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[69] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[70] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
RAM_INST[71] = 32'b000001_11101_00100_0000000000000100; // lw 4 $fp 4
RAM_INST[72] = 32'b000000_00011_00100_00011_00000_000101; // add 3 3 4
RAM_INST[73] = 32'b000010_00011_00010_0000000000000000; // sw 2 3 0
RAM_INST[74] = 32'b000001_11101_00010_0000000000000101; // lw 2 $fp 5
RAM_INST[75] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
RAM_INST[76] = 32'b000001_11101_00100_0000000000000011; // lw 4 $fp 3
RAM_INST[77] = 32'b000000_00011_00100_00011_00000_000101; // add 3 3 4
RAM_INST[78] = 32'b000010_00011_00010_0000000000000000; // sw 2 3 0
RAM_INST[79] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3
RAM_INST[80] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
RAM_INST[81] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
RAM_INST[82] = 32'b001011_00000000000000000000101101; // jump _WhileBegin1_
RAM_INST[83] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit1_
RAM_INST[84] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[85] = 32'b001111_11110_11111_0000000000000000; // push $ra / gcd
RAM_INST[86] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1
RAM_INST[87] = 32'b000101_00000_00011_0000000000000000; // li 3 0
RAM_INST[88] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[89] = 32'b000111_00010_00000_0000000000000110; // beq 2 $zero _ElseBegin1_
RAM_INST[90] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[91] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[92] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[93] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[94] = 32'b001011_00000000000000000001110000; // jump _IfExit1_
RAM_INST[95] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1 / _ElseBegin1_
RAM_INST[96] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
RAM_INST[97] = 32'b000001_11101_00100_0000000000000000; // lw 4 $fp 0
RAM_INST[98] = 32'b000001_11101_00101_0000000000000001; // lw 5 $fp 1
RAM_INST[99] = 32'b000000_00100_00101_00100_00000_001000; // div 4 4 5
RAM_INST[100] = 32'b000001_11101_00101_0000000000000001; // lw 5 $fp 1
RAM_INST[101] = 32'b000000_00100_00101_00100_00000_000111; // mult 4 4 5
RAM_INST[102] = 32'b000000_00011_00100_00011_00000_000110; // sub 3 3 4
RAM_INST[103] = 32'b000011_11101_11101_0000000000000010; // addi $fp $fp 2
RAM_INST[104] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[105] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[106] = 32'b001100_00000000000000000001010101; // jal gcd
RAM_INST[107] = 32'b000100_11101_11101_0000000000000010; // subi $fp $fp 2
RAM_INST[108] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[109] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[110] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[111] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[112] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit1_
RAM_INST[113] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[114] = 32'b001111_11110_11111_0000000000000000; // push $ra / fibonacci
RAM_INST[115] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[116] = 32'b000101_00000_00011_0000000000000000; // li 3 0
RAM_INST[117] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
RAM_INST[118] = 32'b000000_00010_00000_00010_00000_010011; // set 2 2 $zero
RAM_INST[119] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin2_
RAM_INST[120] = 32'b000101_00000_11100_0000000000000000; // li $rv 0
RAM_INST[121] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[122] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[123] = 32'b001011_00000000000000000010011101; // jump _IfExit2_
RAM_INST[124] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin2_
RAM_INST[125] = 32'b000101_00000_00011_0000000000000001; // li 3 1
RAM_INST[126] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[127] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin3_
RAM_INST[128] = 32'b000101_00000_11100_0000000000000001; // li $rv 1
RAM_INST[129] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[130] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[131] = 32'b001011_00000000000000000010011101; // jump _IfExit3_
RAM_INST[132] = 32'b000101_00000_00010_0000000000000000; // li 2 0 / _ElseBegin3_
RAM_INST[133] = 32'b000010_11101_00010_0000000000000001; // sw 2 $fp 1
RAM_INST[134] = 32'b000101_00000_00010_0000000000000001; // li 2 1
RAM_INST[135] = 32'b000010_11101_00010_0000000000000100; // sw 2 $fp 4
RAM_INST[136] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[137] = 32'b000001_11101_00010_0000000000000100; // lw 2 $fp 4 / _WhileBegin2_
RAM_INST[138] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
RAM_INST[139] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[140] = 32'b000111_00010_00000_0000000000001101; // beq 2 $zero _WhileExit2_
RAM_INST[141] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2
RAM_INST[142] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
RAM_INST[143] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2
RAM_INST[144] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[145] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[146] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[147] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3
RAM_INST[148] = 32'b000010_11101_00010_0000000000000001; // sw 2 $fp 1
RAM_INST[149] = 32'b000001_11101_00010_0000000000000100; // lw 2 $fp 4
RAM_INST[150] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
RAM_INST[151] = 32'b000010_11101_00010_0000000000000100; // sw 2 $fp 4
RAM_INST[152] = 32'b001011_00000000000000000010001001; // jump _WhileBegin2_
RAM_INST[153] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _WhileExit2_
RAM_INST[154] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[155] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[156] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[157] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit3_ _IfExit2_
RAM_INST[158] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[159] = 32'b001111_11110_11111_0000000000000000; // push $ra / buscaBinariaInterno
RAM_INST[160] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2
RAM_INST[161] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[162] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[163] = 32'b000101_00000_00011_0000000000000010; // li 3 2
RAM_INST[164] = 32'b000000_00010_00011_00010_00000_001000; // div 2 2 3
RAM_INST[165] = 32'b000010_11101_00010_0000000000000100; // sw 2 $fp 4
RAM_INST[166] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2
RAM_INST[167] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[168] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[169] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin4_
RAM_INST[170] = 32'b000101_00000_11100_0000000000000000; // li $rv 0
RAM_INST[171] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[172] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[173] = 32'b001011_00000000000000000011100100; // jump _IfExit4_
RAM_INST[174] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3 / _ElseBegin4_
RAM_INST[175] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
RAM_INST[176] = 32'b000001_11101_00100_0000000000000100; // lw 4 $fp 4
RAM_INST[177] = 32'b000100_00100_00100_0000000000000001; // subi 4 4 1
RAM_INST[178] = 32'b000000_00011_00100_00011_00000_000101; // add 3 3 4
RAM_INST[179] = 32'b000001_00011_00011_0000000000000000; // lw 3 3 0
RAM_INST[180] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
RAM_INST[181] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin5_
RAM_INST[182] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[183] = 32'b000001_11101_00011_0000000000000100; // lw 3 $fp 4
RAM_INST[184] = 32'b000011_00011_00011_0000000000000001; // addi 3 3 1
RAM_INST[185] = 32'b000001_11101_00100_0000000000000010; // lw 4 $fp 2
RAM_INST[186] = 32'b000001_11101_00101_0000000000000011; // lw 5 $fp 3
RAM_INST[187] = 32'b000011_11101_11101_0000000000000101; // addi $fp $fp 5
RAM_INST[188] = 32'b000010_11101_00101_0000000000000011; // sw 5 $fp 3
RAM_INST[189] = 32'b000010_11101_00100_0000000000000010; // sw 4 $fp 2
RAM_INST[190] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[191] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[192] = 32'b001100_00000000000000000010011111; // jal buscaBinariaInterno
RAM_INST[193] = 32'b000100_11101_11101_0000000000000101; // subi $fp $fp 5
RAM_INST[194] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[195] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[196] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[197] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[198] = 32'b001011_00000000000000000011100100; // jump _IfExit5_
RAM_INST[199] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3 / _ElseBegin5_
RAM_INST[200] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
RAM_INST[201] = 32'b000001_11101_00100_0000000000000100; // lw 4 $fp 4
RAM_INST[202] = 32'b000100_00100_00100_0000000000000001; // subi 4 4 1
RAM_INST[203] = 32'b000000_00011_00100_00011_00000_000101; // add 3 3 4
RAM_INST[204] = 32'b000001_00011_00011_0000000000000000; // lw 3 3 0
RAM_INST[205] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[206] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _ElseBegin6_
RAM_INST[207] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[208] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[209] = 32'b000001_11101_00100_0000000000000100; // lw 4 $fp 4
RAM_INST[210] = 32'b000100_00100_00100_0000000000000001; // subi 4 4 1
RAM_INST[211] = 32'b000001_11101_00101_0000000000000011; // lw 5 $fp 3
RAM_INST[212] = 32'b000011_11101_11101_0000000000000101; // addi $fp $fp 5
RAM_INST[213] = 32'b000010_11101_00101_0000000000000011; // sw 5 $fp 3
RAM_INST[214] = 32'b000010_11101_00100_0000000000000010; // sw 4 $fp 2
RAM_INST[215] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[216] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[217] = 32'b001100_00000000000000000010011111; // jal buscaBinariaInterno
RAM_INST[218] = 32'b000100_11101_11101_0000000000000101; // subi $fp $fp 5
RAM_INST[219] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[220] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[221] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[222] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[223] = 32'b001011_00000000000000000011100100; // jump _IfExit6_
RAM_INST[224] = 32'b000001_11101_00010_0000000000000100; // lw 2 $fp 4 / _ElseBegin6_
RAM_INST[225] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[226] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[227] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[228] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit6_ _IfExit5_ _IfExit4_
RAM_INST[229] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[230] = 32'b001111_11110_11111_0000000000000000; // push $ra / buscaBinaria
RAM_INST[231] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[232] = 32'b000101_00000_00011_0000000000000001; // li 3 1
RAM_INST[233] = 32'b000001_11101_00100_0000000000000001; // lw 4 $fp 1
RAM_INST[234] = 32'b000001_11101_00101_0000000000000010; // lw 5 $fp 2
RAM_INST[235] = 32'b000011_11101_11101_0000000000000011; // addi $fp $fp 3
RAM_INST[236] = 32'b000010_11101_00101_0000000000000011; // sw 5 $fp 3
RAM_INST[237] = 32'b000010_11101_00100_0000000000000010; // sw 4 $fp 2
RAM_INST[238] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[239] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[240] = 32'b001100_00000000000000000010011111; // jal buscaBinariaInterno
RAM_INST[241] = 32'b000100_11101_11101_0000000000000011; // subi $fp $fp 3
RAM_INST[242] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[243] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[244] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[245] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[246] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[247] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[248] = 32'b001111_11110_11111_0000000000000000; // push $ra / fatorial
RAM_INST[249] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[250] = 32'b000101_00000_00011_0000000000000010; // li 3 2
RAM_INST[251] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[252] = 32'b000111_00010_00000_0000000000000101; // beq 2 $zero _ElseBegin7_
RAM_INST[253] = 32'b000101_00000_11100_0000000000000001; // li $rv 1
RAM_INST[254] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[255] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[256] = 32'b001011_00000000000000000100001101; // jump _IfExit7_
RAM_INST[257] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin7_
RAM_INST[258] = 32'b000100_00010_00010_0000000000000001; // subi 2 2 1
RAM_INST[259] = 32'b000011_11101_11101_0000000000000001; // addi $fp $fp 1
RAM_INST[260] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[261] = 32'b001100_00000000000000000011111000; // jal fatorial
RAM_INST[262] = 32'b000100_11101_11101_0000000000000001; // subi $fp $fp 1
RAM_INST[263] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[264] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
RAM_INST[265] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
RAM_INST[266] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[267] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[268] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[269] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit7_
RAM_INST[270] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[271] = 32'b001111_11110_11111_0000000000000000; // push $ra / calculadora
RAM_INST[272] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2
RAM_INST[273] = 32'b000101_00000_00011_0000000000000001; // li 3 1
RAM_INST[274] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[275] = 32'b000111_00010_00000_0000000000001000; // beq 2 $zero _ElseBegin8_
RAM_INST[276] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[277] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[278] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[279] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[280] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[281] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[282] = 32'b001011_00000000000000000101011011; // jump _IfExit8_
RAM_INST[283] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _ElseBegin8_
RAM_INST[284] = 32'b000101_00000_00011_0000000000000010; // li 3 2
RAM_INST[285] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[286] = 32'b000111_00010_00000_0000000000001000; // beq 2 $zero _ElseBegin9_
RAM_INST[287] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[288] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[289] = 32'b000000_00010_00011_00010_00000_000110; // sub 2 2 3
RAM_INST[290] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[291] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[292] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[293] = 32'b001011_00000000000000000101011011; // jump _IfExit9_
RAM_INST[294] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _ElseBegin9_
RAM_INST[295] = 32'b000101_00000_00011_0000000000000011; // li 3 3
RAM_INST[296] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[297] = 32'b000111_00010_00000_0000000000001000; // beq 2 $zero _ElseBegin10_
RAM_INST[298] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[299] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[300] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
RAM_INST[301] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[302] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[303] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[304] = 32'b001011_00000000000000000101011011; // jump _IfExit10_
RAM_INST[305] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _ElseBegin10_
RAM_INST[306] = 32'b000101_00000_00011_0000000000000100; // li 3 4
RAM_INST[307] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[308] = 32'b000111_00010_00000_0000000000001000; // beq 2 $zero _ElseBegin11_
RAM_INST[309] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[310] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[311] = 32'b000000_00010_00011_00010_00000_001000; // div 2 2 3
RAM_INST[312] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[313] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[314] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[315] = 32'b001011_00000000000000000101011011; // jump _IfExit11_
RAM_INST[316] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _ElseBegin11_
RAM_INST[317] = 32'b000101_00000_00011_0000000000000101; // li 3 5
RAM_INST[318] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[319] = 32'b000111_00010_00000_0000000000001100; // beq 2 $zero _ElseBegin12_
RAM_INST[320] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[321] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
RAM_INST[322] = 32'b000001_11101_00100_0000000000000001; // lw 4 $fp 1
RAM_INST[323] = 32'b000000_00011_00100_00011_00000_001000; // div 3 3 4
RAM_INST[324] = 32'b000001_11101_00100_0000000000000001; // lw 4 $fp 1
RAM_INST[325] = 32'b000000_00011_00100_00011_00000_000111; // mult 3 3 4
RAM_INST[326] = 32'b000000_00010_00011_00010_00000_000110; // sub 2 2 3
RAM_INST[327] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[328] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[329] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[330] = 32'b001011_00000000000000000101011011; // jump _IfExit12_
RAM_INST[331] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _ElseBegin12_
RAM_INST[332] = 32'b000101_00000_00011_0000000000000110; // li 3 6
RAM_INST[333] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[334] = 32'b000111_00010_00000_0000000000001010; // beq 2 $zero _ElseBegin13_
RAM_INST[335] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[336] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[337] = 32'b000000_00010_00011_00010_00000_000111; // mult 2 2 3
RAM_INST[338] = 32'b000101_00000_00011_0000000001100100; // li 3 100
RAM_INST[339] = 32'b000000_00010_00011_00010_00000_001000; // div 2 2 3
RAM_INST[340] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[341] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[342] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[343] = 32'b001011_00000000000000000101011011; // jump _IfExit13_
RAM_INST[344] = 32'b000101_00000_11100_0000000000000000; // li $rv 0 / _ElseBegin13_
RAM_INST[345] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[346] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[347] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _IfExit13_ _IfExit12_ _IfExit11_ _IfExit10_ _IfExit9_ _IfExit8_
RAM_INST[348] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[349] = 32'b001111_11110_11111_0000000000000000; // push $ra / mediaVector
RAM_INST[350] = 32'b000101_00000_00010_0000000000000000; // li 2 0
RAM_INST[351] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[352] = 32'b000101_00000_00010_0000000000000000; // li 2 0
RAM_INST[353] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
RAM_INST[354] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _WhileBegin3_
RAM_INST[355] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[356] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[357] = 32'b000111_00010_00000_0000000000001100; // beq 2 $zero _WhileExit3_
RAM_INST[358] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3
RAM_INST[359] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
RAM_INST[360] = 32'b000001_11101_00100_0000000000000010; // lw 4 $fp 2
RAM_INST[361] = 32'b000000_00011_00100_00011_00000_000101; // add 3 3 4
RAM_INST[362] = 32'b000001_00011_00011_0000000000000000; // lw 3 3 0
RAM_INST[363] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[364] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
RAM_INST[365] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2
RAM_INST[366] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
RAM_INST[367] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[368] = 32'b001011_00000000000000000101100010; // jump _WhileBegin3_
RAM_INST[369] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3 / _WhileExit3_
RAM_INST[370] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[371] = 32'b000000_00010_00011_00010_00000_001000; // div 2 2 3
RAM_INST[372] = 32'b000000_00010_11100_00000_00000_010000; // move $rv 2
RAM_INST[373] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[374] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[375] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[376] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[377] = 32'b001111_11110_11111_0000000000000000; // push $ra / extremosVector
RAM_INST[378] = 32'b000101_00000_00010_0000000000000001; // li 2 1
RAM_INST[379] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[380] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[381] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[382] = 32'b000010_11101_00010_0000000000000100; // sw 2 $fp 4
RAM_INST[383] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
RAM_INST[384] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _WhileBegin4_
RAM_INST[385] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[386] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[387] = 32'b000111_00010_00000_0000000000011110; // beq 2 $zero _WhileExit4_
RAM_INST[388] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[389] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
RAM_INST[390] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[391] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[392] = 32'b000001_11101_00011_0000000000000011; // lw 3 $fp 3
RAM_INST[393] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[394] = 32'b000111_00010_00000_0000000000000111; // beq 2 $zero _ElseBegin14_
RAM_INST[395] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[396] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
RAM_INST[397] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[398] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[399] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
RAM_INST[400] = 32'b001011_00000000000000000110011101; // jump _IfExit14_
RAM_INST[401] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin14_
RAM_INST[402] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
RAM_INST[403] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[404] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[405] = 32'b000001_11101_00011_0000000000000100; // lw 3 $fp 4
RAM_INST[406] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
RAM_INST[407] = 32'b000111_00010_00000_0000000000000110; // beq 2 $zero _IfExit15_
RAM_INST[408] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[409] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
RAM_INST[410] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[411] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[412] = 32'b000010_11101_00010_0000000000000100; // sw 2 $fp 4
RAM_INST[413] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _IfExit15_ _IfExit14_
RAM_INST[414] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
RAM_INST[415] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[416] = 32'b001011_00000000000000000110000000; // jump _WhileBegin4_
RAM_INST[417] = 32'b000001_11101_00010_0000000000000011; // lw 2 $fp 3 / _WhileExit4_
RAM_INST[418] = 32'b001010_00010_00000_0000000000000000; // out 2
RAM_INST[419] = 32'b000001_11101_00010_0000000000000100; // lw 2 $fp 4
RAM_INST[420] = 32'b001010_00010_00000_0000000000000000; // out 2
RAM_INST[421] = 32'b010000_11110_11111_0000000000000000; // pop $ra
RAM_INST[422] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[423] = 32'b001111_11110_11111_0000000000000000; // push $ra / inputVector
RAM_INST[424] = 32'b000101_00000_00010_0000000000000000; // li 2 0
RAM_INST[425] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[426] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _WhileBegin5_
RAM_INST[427] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[428] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[429] = 32'b000111_00010_00000_0000000000001010; // beq 2 $zero _WhileExit5_
RAM_INST[430] = 32'b001001_00000_00010_0000000000000000; // in 2
RAM_INST[431] = 32'b000001_11101_00011_0000000000000000; // lw 3 $fp 0
RAM_INST[432] = 32'b000001_11101_00100_0000000000000010; // lw 4 $fp 2
RAM_INST[433] = 32'b000000_00011_00100_00011_00000_000101; // add 3 3 4
RAM_INST[434] = 32'b000010_00011_00010_0000000000000000; // sw 2 3 0
RAM_INST[435] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2
RAM_INST[436] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
RAM_INST[437] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[438] = 32'b001011_00000000000000000110101010; // jump _WhileBegin5_
RAM_INST[439] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit5_
RAM_INST[440] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[441] = 32'b001111_11110_11111_0000000000000000; // push $ra / outputVector
RAM_INST[442] = 32'b000101_00000_00010_0000000000000000; // li 2 0
RAM_INST[443] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[444] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2 / _WhileBegin6_
RAM_INST[445] = 32'b000001_11101_00011_0000000000000001; // lw 3 $fp 1
RAM_INST[446] = 32'b000000_00010_00011_00010_00000_010001; // slt 2 2 3
RAM_INST[447] = 32'b000111_00010_00000_0000000000001010; // beq 2 $zero _WhileExit6_
RAM_INST[448] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[449] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
RAM_INST[450] = 32'b000000_00010_00011_00010_00000_000101; // add 2 2 3
RAM_INST[451] = 32'b000001_00010_00010_0000000000000000; // lw 2 2 0
RAM_INST[452] = 32'b001010_00010_00000_0000000000000000; // out 2
RAM_INST[453] = 32'b000001_11101_00010_0000000000000010; // lw 2 $fp 2
RAM_INST[454] = 32'b000011_00010_00010_0000000000000001; // addi 2 2 1
RAM_INST[455] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[456] = 32'b001011_00000000000000000110111100; // jump _WhileBegin6_
RAM_INST[457] = 32'b010000_11110_11111_0000000000000000; // pop $ra / _WhileExit6_
RAM_INST[458] = 32'b000000_11111_00000_00000_00000_010100; // jr $ra
RAM_INST[459] = 32'b001001_00000_00010_0000000000000000; // in 2 / main
RAM_INST[460] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[461] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _WhileBegin7_
RAM_INST[462] = 32'b000101_00000_00011_0000000000000000; // li 3 0
RAM_INST[463] = 32'b000000_00010_00011_00010_00000_010010; // sgt 2 2 3
RAM_INST[464] = 32'b000111_00010_00000_0000000010010101; // beq 2 $zero _WhileExit7_
RAM_INST[465] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0
RAM_INST[466] = 32'b000101_00000_00011_0000000000000001; // li 3 1
RAM_INST[467] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[468] = 32'b000111_00010_00000_0000000000001001; // beq 2 $zero _ElseBegin16_
RAM_INST[469] = 32'b000011_11011_00010_0000000000000000; // addi 2 $global 0
RAM_INST[470] = 32'b000101_00000_00011_0000000000001010; // li 3 10
RAM_INST[471] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
RAM_INST[472] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[473] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[474] = 32'b001100_00000000000000000110100111; // jal inputVector
RAM_INST[475] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
RAM_INST[476] = 32'b001011_00000000000000001001100010; // jump _IfExit16_
RAM_INST[477] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin16_
RAM_INST[478] = 32'b000101_00000_00011_0000000000000010; // li 3 2
RAM_INST[479] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[480] = 32'b000111_00010_00000_0000000000001001; // beq 2 $zero _ElseBegin17_
RAM_INST[481] = 32'b000011_11011_00010_0000000000000000; // addi 2 $global 0
RAM_INST[482] = 32'b000101_00000_00011_0000000000001010; // li 3 10
RAM_INST[483] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
RAM_INST[484] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[485] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[486] = 32'b001100_00000000000000000110111001; // jal outputVector
RAM_INST[487] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
RAM_INST[488] = 32'b001011_00000000000000001001100010; // jump _IfExit17_
RAM_INST[489] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin17_
RAM_INST[490] = 32'b000101_00000_00011_0000000000000011; // li 3 3
RAM_INST[491] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[492] = 32'b000111_00010_00000_0000000000001011; // beq 2 $zero _ElseBegin18_
RAM_INST[493] = 32'b000011_11011_00010_0000000000000000; // addi 2 $global 0
RAM_INST[494] = 32'b000101_00000_00011_0000000000000000; // li 3 0
RAM_INST[495] = 32'b000101_00000_00100_0000000000001010; // li 4 10
RAM_INST[496] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
RAM_INST[497] = 32'b000010_11101_00100_0000000000000010; // sw 4 $fp 2
RAM_INST[498] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[499] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[500] = 32'b001100_00000000000000000000101010; // jal sort
RAM_INST[501] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
RAM_INST[502] = 32'b001011_00000000000000001001100010; // jump _IfExit18_
RAM_INST[503] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin18_
RAM_INST[504] = 32'b000101_00000_00011_0000000000000100; // li 3 4
RAM_INST[505] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[506] = 32'b000111_00010_00000_0000000000001011; // beq 2 $zero _ElseBegin19_
RAM_INST[507] = 32'b000011_11011_00010_0000000000000000; // addi 2 $global 0
RAM_INST[508] = 32'b000101_00000_00011_0000000000001010; // li 3 10
RAM_INST[509] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
RAM_INST[510] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[511] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[512] = 32'b001100_00000000000000000101011101; // jal mediaVector
RAM_INST[513] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
RAM_INST[514] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[515] = 32'b001010_00010_00000_0000000000000000; // out 2
RAM_INST[516] = 32'b001011_00000000000000001001100010; // jump _IfExit19_
RAM_INST[517] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin19_
RAM_INST[518] = 32'b000101_00000_00011_0000000000000101; // li 3 5
RAM_INST[519] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[520] = 32'b000111_00010_00000_0000000000001001; // beq 2 $zero _ElseBegin20_
RAM_INST[521] = 32'b000011_11011_00010_0000000000000000; // addi 2 $global 0
RAM_INST[522] = 32'b000101_00000_00011_0000000000001010; // li 3 10
RAM_INST[523] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
RAM_INST[524] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[525] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[526] = 32'b001100_00000000000000000101111001; // jal extremosVector
RAM_INST[527] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
RAM_INST[528] = 32'b001011_00000000000000001001100010; // jump _IfExit20_
RAM_INST[529] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin20_
RAM_INST[530] = 32'b000101_00000_00011_0000000000000110; // li 3 6
RAM_INST[531] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[532] = 32'b000111_00010_00000_0000000000001111; // beq 2 $zero _ElseBegin21_
RAM_INST[533] = 32'b001001_00000_00010_0000000000000000; // in 2
RAM_INST[534] = 32'b000010_11101_00010_0000000000000001; // sw 2 $fp 1
RAM_INST[535] = 32'b000011_11011_00010_0000000000000000; // addi 2 $global 0
RAM_INST[536] = 32'b000101_00000_00011_0000000000001010; // li 3 10
RAM_INST[537] = 32'b000001_11101_00100_0000000000000001; // lw 4 $fp 1
RAM_INST[538] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
RAM_INST[539] = 32'b000010_11101_00100_0000000000000010; // sw 4 $fp 2
RAM_INST[540] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[541] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[542] = 32'b001100_00000000000000000011100110; // jal buscaBinaria
RAM_INST[543] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
RAM_INST[544] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[545] = 32'b001010_00010_00000_0000000000000000; // out 2
RAM_INST[546] = 32'b001011_00000000000000001001100010; // jump _IfExit21_
RAM_INST[547] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin21_
RAM_INST[548] = 32'b000101_00000_00011_0000000000000111; // li 3 7
RAM_INST[549] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[550] = 32'b000111_00010_00000_0000000000001111; // beq 2 $zero _ElseBegin22_
RAM_INST[551] = 32'b001001_00000_00010_0000000000000000; // in 2
RAM_INST[552] = 32'b000010_11101_00010_0000000000000001; // sw 2 $fp 1
RAM_INST[553] = 32'b001001_00000_00010_0000000000000000; // in 2
RAM_INST[554] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[555] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1
RAM_INST[556] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
RAM_INST[557] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
RAM_INST[558] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[559] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[560] = 32'b001100_00000000000000000001010101; // jal gcd
RAM_INST[561] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
RAM_INST[562] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[563] = 32'b001010_00010_00000_0000000000000000; // out 2
RAM_INST[564] = 32'b001011_00000000000000001001100010; // jump _IfExit22_
RAM_INST[565] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin22_
RAM_INST[566] = 32'b000101_00000_00011_0000000000001000; // li 3 8
RAM_INST[567] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[568] = 32'b000111_00010_00000_0000000000001001; // beq 2 $zero _ElseBegin23_
RAM_INST[569] = 32'b001001_00000_00010_0000000000000000; // in 2
RAM_INST[570] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
RAM_INST[571] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[572] = 32'b001100_00000000000000000001110010; // jal fibonacci
RAM_INST[573] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
RAM_INST[574] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[575] = 32'b001010_00010_00000_0000000000000000; // out 2
RAM_INST[576] = 32'b001011_00000000000000001001100010; // jump _IfExit23_
RAM_INST[577] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin23_
RAM_INST[578] = 32'b000101_00000_00011_0000000000001001; // li 3 9
RAM_INST[579] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[580] = 32'b000111_00010_00000_0000000000001001; // beq 2 $zero _ElseBegin24_
RAM_INST[581] = 32'b001001_00000_00010_0000000000000000; // in 2
RAM_INST[582] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
RAM_INST[583] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[584] = 32'b001100_00000000000000000011111000; // jal fatorial
RAM_INST[585] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
RAM_INST[586] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[587] = 32'b001010_00010_00000_0000000000000000; // out 2
RAM_INST[588] = 32'b001011_00000000000000001001100010; // jump _IfExit24_
RAM_INST[589] = 32'b000001_11101_00010_0000000000000000; // lw 2 $fp 0 / _ElseBegin24_
RAM_INST[590] = 32'b000101_00000_00011_0000000000001010; // li 3 10
RAM_INST[591] = 32'b000000_00010_00011_00010_00000_010011; // set 2 2 3
RAM_INST[592] = 32'b000111_00010_00000_0000000000010010; // beq 2 $zero _IfExit25_
RAM_INST[593] = 32'b001001_00000_00010_0000000000000000; // in 2
RAM_INST[594] = 32'b000010_11101_00010_0000000000000001; // sw 2 $fp 1
RAM_INST[595] = 32'b001001_00000_00010_0000000000000000; // in 2
RAM_INST[596] = 32'b000010_11101_00010_0000000000000010; // sw 2 $fp 2
RAM_INST[597] = 32'b001001_00000_00010_0000000000000000; // in 2
RAM_INST[598] = 32'b000010_11101_00010_0000000000000011; // sw 2 $fp 3
RAM_INST[599] = 32'b000001_11101_00010_0000000000000001; // lw 2 $fp 1
RAM_INST[600] = 32'b000001_11101_00011_0000000000000010; // lw 3 $fp 2
RAM_INST[601] = 32'b000001_11101_00100_0000000000000011; // lw 4 $fp 3
RAM_INST[602] = 32'b000011_11101_11101_0000000000000100; // addi $fp $fp 4
RAM_INST[603] = 32'b000010_11101_00100_0000000000000010; // sw 4 $fp 2
RAM_INST[604] = 32'b000010_11101_00011_0000000000000001; // sw 3 $fp 1
RAM_INST[605] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[606] = 32'b001100_00000000000000000100001111; // jal calculadora
RAM_INST[607] = 32'b000100_11101_11101_0000000000000100; // subi $fp $fp 4
RAM_INST[608] = 32'b000000_11100_00010_00000_00000_010000; // move 2 $rv
RAM_INST[609] = 32'b001010_00010_00000_0000000000000000; // out 2
RAM_INST[610] = 32'b001001_00000_00010_0000000000000000; // in 2 / _IfExit25_ _IfExit24_ _IfExit23_ _IfExit22_ _IfExit21_ _IfExit20_ _IfExit19_ _IfExit18_ _IfExit17_ _IfExit16_
RAM_INST[611] = 32'b000010_11101_00010_0000000000000000; // sw 2 $fp 0
RAM_INST[612] = 32'b001011_00000000000000000111001101; // jump _WhileBegin7_
RAM_INST[613] = 32'b11111111111111111111111111111111; // halt / _halt_ _WhileExit7_
*/
			
		end

		
	end
	
	always @ (posedge read_clock)
	begin
		
		out <= RAM_INST[memAddress];
		
	end
	
	
	
endmodule

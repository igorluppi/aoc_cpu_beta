module freq_div (clk, clk_out);
	input clk;
	output reg clk_out = 0;
	reg [13:0] estado = 0;

	always@(posedge clk)
		begin
			/*case(estado)
				0: estado = 1;
1: estado = 2;
2: estado = 3;
3: estado = 4;
4: estado = 5;
5: estado = 6;
6: estado = 7;
7: estado = 8;
8: estado = 9;
9: estado = 10;
10: estado = 11;
11: estado = 12;
12: estado = 13;
13: estado = 14;
14: estado = 15;
15: estado = 16;
16: estado = 17;
17: estado = 18;
18: estado = 19;
19: estado = 20;
20: estado = 21;
21: estado = 22;
22: estado = 23;
23: estado = 24;
24: estado = 25;
25: estado = 26;
26: estado = 27;
27: estado = 28;
28: estado = 29;
29: estado = 30;
30: estado = 31;
31: estado = 32;
32: estado = 33;
33: estado = 34;
34: estado = 35;
35: estado = 36;
36: estado = 37;
37: estado = 38;
38: estado = 39;
39: estado = 40;
40: estado = 41;
41: estado = 42;
42: estado = 43;
43: estado = 44;
44: estado = 45;
45: estado = 46;
46: estado = 47;
47: estado = 48;
48: estado = 49;
49: estado = 50;
50: estado = 51;
51: estado = 52;
52: estado = 53;
53: estado = 54;
54: estado = 55;
55: estado = 56;
56: estado = 57;
57: estado = 58;
58: estado = 59;
59: estado = 60;
60: estado = 61;
61: estado = 62;
62: estado = 63;
63: estado = 64;
64: estado = 65;
65: estado = 66;
66: estado = 67;
67: estado = 68;
68: estado = 69;
69: estado = 70;
70: estado = 71;
71: estado = 72;
72: estado = 73;
73: estado = 74;
74: estado = 75;
75: estado = 76;
76: estado = 77;
77: estado = 78;
78: estado = 79;
79: estado = 80;
80: estado = 81;
81: estado = 82;
82: estado = 83;
83: estado = 84;
84: estado = 85;
85: estado = 86;
86: estado = 87;
87: estado = 88;
88: estado = 89;
89: estado = 90;
90: estado = 91;
91: estado = 92;
92: estado = 93;
93: estado = 94;
94: estado = 95;
95: estado = 96;
96: estado = 97;
97: estado = 98;
98: estado = 99;
99: estado = 100;
100: estado = 101;
101: estado = 102;
102: estado = 103;
103: estado = 104;
104: estado = 105;
105: estado = 106;
106: estado = 107;
107: estado = 108;
108: estado = 109;
109: estado = 110;
110: estado = 111;
111: estado = 112;
112: estado = 113;
113: estado = 114;
114: estado = 115;
115: estado = 116;
116: estado = 117;
117: estado = 118;
118: estado = 119;
119: estado = 120;
120: estado = 121;
121: estado = 122;
122: estado = 123;
123: estado = 124;
124: estado = 125;
125: estado = 126;
126: estado = 127;
127: estado = 128;
128: estado = 129;
129: estado = 130;
130: estado = 131;
131: estado = 132;
132: estado = 133;
133: estado = 134;
134: estado = 135;
135: estado = 136;
136: estado = 137;
137: estado = 138;
138: estado = 139;
139: estado = 140;
140: estado = 141;
141: estado = 142;
142: estado = 143;
143: estado = 144;
144: estado = 145;
145: estado = 146;
146: estado = 147;
147: estado = 148;
148: estado = 149;
149: estado = 150;
150: estado = 151;
151: estado = 152;
152: estado = 153;
153: estado = 154;
154: estado = 155;
155: estado = 156;
156: estado = 157;
157: estado = 158;
158: estado = 159;
159: estado = 160;
160: estado = 161;
161: estado = 162;
162: estado = 163;
163: estado = 164;
164: estado = 165;
165: estado = 166;
166: estado = 167;
167: estado = 168;
168: estado = 169;
169: estado = 170;
170: estado = 171;
171: estado = 172;
172: estado = 173;
173: estado = 174;
174: estado = 175;
175: estado = 176;
176: estado = 177;
177: estado = 178;
178: estado = 179;
179: estado = 180;
180: estado = 181;
181: estado = 182;
182: estado = 183;
183: estado = 184;
184: estado = 185;
185: estado = 186;
186: estado = 187;
187: estado = 188;
188: estado = 189;
189: estado = 190;
190: estado = 191;
191: estado = 192;
192: estado = 193;
193: estado = 194;
194: estado = 195;
195: estado = 196;
196: estado = 197;
197: estado = 198;
198: estado = 199;
199: estado = 200;
200: estado = 201;
201: estado = 202;
202: estado = 203;
203: estado = 204;
204: estado = 205;
205: estado = 206;
206: estado = 207;
207: estado = 208;
208: estado = 209;
209: estado = 210;
210: estado = 211;
211: estado = 212;
212: estado = 213;
213: estado = 214;
214: estado = 215;
215: estado = 216;
216: estado = 217;
217: estado = 218;
218: estado = 219;
219: estado = 220;
220: estado = 221;
221: estado = 222;
222: estado = 223;
223: estado = 224;
224: estado = 225;
225: estado = 226;
226: estado = 227;
227: estado = 228;
228: estado = 229;
229: estado = 230;
230: estado = 231;
231: estado = 232;
232: estado = 233;
233: estado = 234;
234: estado = 235;
235: estado = 236;
236: estado = 237;
237: estado = 238;
238: estado = 239;
239: estado = 240;
240: estado = 241;
241: estado = 242;
242: estado = 243;
243: estado = 244;
244: estado = 245;
245: estado = 246;
246: estado = 247;
247: estado = 248;
248: estado = 249;
249: estado = 250;
250: estado = 251;
251: estado = 252;
252: estado = 253;
253: estado = 254;
254: estado = 255;
255: estado = 256;
256: estado = 257;
257: estado = 258;
258: estado = 259;
259: estado = 260;
260: estado = 261;
261: estado = 262;
262: estado = 263;
263: estado = 264;
264: estado = 265;
265: estado = 266;
266: estado = 267;
267: estado = 268;
268: estado = 269;
269: estado = 270;
270: estado = 271;
271: estado = 272;
272: estado = 273;
273: estado = 274;
274: estado = 275;
275: estado = 276;
276: estado = 277;
277: estado = 278;
278: estado = 279;
279: estado = 280;
280: estado = 281;
281: estado = 282;
282: estado = 283;
283: estado = 284;
284: estado = 285;
285: estado = 286;
286: estado = 287;
287: estado = 288;
288: estado = 289;
289: estado = 290;
290: estado = 291;
291: estado = 292;
292: estado = 293;
293: estado = 294;
294: estado = 295;
295: estado = 296;
296: estado = 297;
297: estado = 298;
298: estado = 299;
299: estado = 300;
300: estado = 301;
301: estado = 302;
302: estado = 303;
303: estado = 304;
304: estado = 305;
305: estado = 306;
306: estado = 307;
307: estado = 308;
308: estado = 309;
309: estado = 310;
310: estado = 311;
311: estado = 312;
312: estado = 313;
313: estado = 314;
314: estado = 315;
315: estado = 316;
316: estado = 317;
317: estado = 318;
318: estado = 319;
319: estado = 320;
320: estado = 321;
321: estado = 322;
322: estado = 323;
323: estado = 324;
324: estado = 325;
325: estado = 326;
326: estado = 327;
327: estado = 328;
328: estado = 329;
329: estado = 330;
330: estado = 331;
331: estado = 332;
332: estado = 333;
333: estado = 334;
334: estado = 335;
335: estado = 336;
336: estado = 337;
337: estado = 338;
338: estado = 339;
339: estado = 340;
340: estado = 341;
341: estado = 342;
342: estado = 343;
343: estado = 344;
344: estado = 345;
345: estado = 346;
346: estado = 347;
347: estado = 348;
348: estado = 349;
349: estado = 350;
350: estado = 351;
351: estado = 352;
352: estado = 353;
353: estado = 354;
354: estado = 355;
355: estado = 356;
356: estado = 357;
357: estado = 358;
358: estado = 359;
359: estado = 360;
360: estado = 361;
361: estado = 362;
362: estado = 363;
363: estado = 364;
364: estado = 365;
365: estado = 366;
366: estado = 367;
367: estado = 368;
368: estado = 369;
369: estado = 370;
370: estado = 371;
371: estado = 372;
372: estado = 373;
373: estado = 374;
374: estado = 375;
375: estado = 376;
376: estado = 377;
377: estado = 378;
378: estado = 379;
379: estado = 380;
380: estado = 381;
381: estado = 382;
382: estado = 383;
383: estado = 384;
384: estado = 385;
385: estado = 386;
386: estado = 387;
387: estado = 388;
388: estado = 389;
389: estado = 390;
390: estado = 391;
391: estado = 392;
392: estado = 393;
393: estado = 394;
394: estado = 395;
395: estado = 396;
396: estado = 397;
397: estado = 398;
398: estado = 399;
399: estado = 400;
400: estado = 401;
401: estado = 402;
402: estado = 403;
403: estado = 404;
404: estado = 405;
405: estado = 406;
406: estado = 407;
407: estado = 408;
408: estado = 409;
409: estado = 410;
410: estado = 411;
411: estado = 412;
412: estado = 413;
413: estado = 414;
414: estado = 415;
415: estado = 416;
416: estado = 417;
417: estado = 418;
418: estado = 419;
419: estado = 420;
420: estado = 421;
421: estado = 422;
422: estado = 423;
423: estado = 424;
424: estado = 425;
425: estado = 426;
426: estado = 427;
427: estado = 428;
428: estado = 429;
429: estado = 430;
430: estado = 431;
431: estado = 432;
432: estado = 433;
433: estado = 434;
434: estado = 435;
435: estado = 436;
436: estado = 437;
437: estado = 438;
438: estado = 439;
439: estado = 440;
440: estado = 441;
441: estado = 442;
442: estado = 443;
443: estado = 444;
444: estado = 445;
445: estado = 446;
446: estado = 447;
447: estado = 448;
448: estado = 449;
449: estado = 450;
450: estado = 451;
451: estado = 452;
452: estado = 453;
453: estado = 454;
454: estado = 455;
455: estado = 456;
456: estado = 457;
457: estado = 458;
458: estado = 459;
459: estado = 460;
460: estado = 461;
461: estado = 462;
462: estado = 463;
463: estado = 464;
464: estado = 465;
465: estado = 466;
466: estado = 467;
467: estado = 468;
468: estado = 469;
469: estado = 470;
470: estado = 471;
471: estado = 472;
472: estado = 473;
473: estado = 474;
474: estado = 475;
475: estado = 476;
476: estado = 477;
477: estado = 478;
478: estado = 479;
479: estado = 480;
480: estado = 481;
481: estado = 482;
482: estado = 483;
483: estado = 484;
484: estado = 485;
485: estado = 486;
486: estado = 487;
487: estado = 488;
488: estado = 489;
489: estado = 490;
490: estado = 491;
491: estado = 492;
492: estado = 493;
493: estado = 494;
494: estado = 495;
495: estado = 496;
496: estado = 497;
497: estado = 498;
498: estado = 499;
499: estado = 500;
500: estado = 501;
501: estado = 502;
502: estado = 503;
503: estado = 504;
504: estado = 505;
505: estado = 506;
506: estado = 507;
507: estado = 508;
508: estado = 509;
509: estado = 510;
510: estado = 511;
511: estado = 512;
512: estado = 513;
513: estado = 514;
514: estado = 515;
515: estado = 516;
516: estado = 517;
517: estado = 518;
518: estado = 519;
519: estado = 520;
520: estado = 521;
521: estado = 522;
522: estado = 523;
523: estado = 524;
524: estado = 525;
525: estado = 526;
526: estado = 527;
527: estado = 528;
528: estado = 529;
529: estado = 530;
530: estado = 531;
531: estado = 532;
532: estado = 533;
533: estado = 534;
534: estado = 535;
535: estado = 536;
536: estado = 537;
537: estado = 538;
538: estado = 539;
539: estado = 540;
540: estado = 541;
541: estado = 542;
542: estado = 543;
543: estado = 544;
544: estado = 545;
545: estado = 546;
546: estado = 547;
547: estado = 548;
548: estado = 549;
549: estado = 550;
550: estado = 551;
551: estado = 552;
552: estado = 553;
553: estado = 554;
554: estado = 555;
555: estado = 556;
556: estado = 557;
557: estado = 558;
558: estado = 559;
559: estado = 560;
560: estado = 561;
561: estado = 562;
562: estado = 563;
563: estado = 564;
564: estado = 565;
565: estado = 566;
566: estado = 567;
567: estado = 568;
568: estado = 569;
569: estado = 570;
570: estado = 571;
571: estado = 572;
572: estado = 573;
573: estado = 574;
574: estado = 575;
575: estado = 576;
576: estado = 577;
577: estado = 578;
578: estado = 579;
579: estado = 580;
580: estado = 581;
581: estado = 582;
582: estado = 583;
583: estado = 584;
584: estado = 585;
585: estado = 586;
586: estado = 587;
587: estado = 588;
588: estado = 589;
589: estado = 590;
590: estado = 591;
591: estado = 592;
592: estado = 593;
593: estado = 594;
594: estado = 595;
595: estado = 596;
596: estado = 597;
597: estado = 598;
598: estado = 599;
599: estado = 600;
600: estado = 601;
601: estado = 602;
602: estado = 603;
603: estado = 604;
604: estado = 605;
605: estado = 606;
606: estado = 607;
607: estado = 608;
608: estado = 609;
609: estado = 610;
610: estado = 611;
611: estado = 612;
612: estado = 613;
613: estado = 614;
614: estado = 615;
615: estado = 616;
616: estado = 617;
617: estado = 618;
618: estado = 619;
619: estado = 620;
620: estado = 621;
621: estado = 622;
622: estado = 623;
623: estado = 624;
624: estado = 625;
625: estado = 626;
626: estado = 627;
627: estado = 628;
628: estado = 629;
629: estado = 630;
630: estado = 631;
631: estado = 632;
632: estado = 633;
633: estado = 634;
634: estado = 635;
635: estado = 636;
636: estado = 637;
637: estado = 638;
638: estado = 639;
639: estado = 640;
640: estado = 641;
641: estado = 642;
642: estado = 643;
643: estado = 644;
644: estado = 645;
645: estado = 646;
646: estado = 647;
647: estado = 648;
648: estado = 649;
649: estado = 650;
650: estado = 651;
651: estado = 652;
652: estado = 653;
653: estado = 654;
654: estado = 655;
655: estado = 656;
656: estado = 657;
657: estado = 658;
658: estado = 659;
659: estado = 660;
660: estado = 661;
661: estado = 662;
662: estado = 663;
663: estado = 664;
664: estado = 665;
665: estado = 666;
666: estado = 667;
667: estado = 668;
668: estado = 669;
669: estado = 670;
670: estado = 671;
671: estado = 672;
672: estado = 673;
673: estado = 674;
674: estado = 675;
675: estado = 676;
676: estado = 677;
677: estado = 678;
678: estado = 679;
679: estado = 680;
680: estado = 681;
681: estado = 682;
682: estado = 683;
683: estado = 684;
684: estado = 685;
685: estado = 686;
686: estado = 687;
687: estado = 688;
688: estado = 689;
689: estado = 690;
690: estado = 691;
691: estado = 692;
692: estado = 693;
693: estado = 694;
694: estado = 695;
695: estado = 696;
696: estado = 697;
697: estado = 698;
698: estado = 699;
699: estado = 700;
700: estado = 701;
701: estado = 702;
702: estado = 703;
703: estado = 704;
704: estado = 705;
705: estado = 706;
706: estado = 707;
707: estado = 708;
708: estado = 709;
709: estado = 710;
710: estado = 711;
711: estado = 712;
712: estado = 713;
713: estado = 714;
714: estado = 715;
715: estado = 716;
716: estado = 717;
717: estado = 718;
718: estado = 719;
719: estado = 720;
720: estado = 721;
721: estado = 722;
722: estado = 723;
723: estado = 724;
724: estado = 725;
725: estado = 726;
726: estado = 727;
727: estado = 728;
728: estado = 729;
729: estado = 730;
730: estado = 731;
731: estado = 732;
732: estado = 733;
733: estado = 734;
734: estado = 735;
735: estado = 736;
736: estado = 737;
737: estado = 738;
738: estado = 739;
739: estado = 740;
740: estado = 741;
741: estado = 742;
742: estado = 743;
743: estado = 744;
744: estado = 745;
745: estado = 746;
746: estado = 747;
747: estado = 748;
748: estado = 749;
749: estado = 750;
750: estado = 751;
751: estado = 752;
752: estado = 753;
753: estado = 754;
754: estado = 755;
755: estado = 756;
756: estado = 757;
757: estado = 758;
758: estado = 759;
759: estado = 760;
760: estado = 761;
761: estado = 762;
762: estado = 763;
763: estado = 764;
764: estado = 765;
765: estado = 766;
766: estado = 767;
767: estado = 768;
768: estado = 769;
769: estado = 770;
770: estado = 771;
771: estado = 772;
772: estado = 773;
773: estado = 774;
774: estado = 775;
775: estado = 776;
776: estado = 777;
777: estado = 778;
778: estado = 779;
779: estado = 780;
780: estado = 781;
781: estado = 782;
782: estado = 783;
783: estado = 784;
784: estado = 785;
785: estado = 786;
786: estado = 787;
787: estado = 788;
788: estado = 789;
789: estado = 790;
790: estado = 791;
791: estado = 792;
792: estado = 793;
793: estado = 794;
794: estado = 795;
795: estado = 796;
796: estado = 797;
797: estado = 798;
798: estado = 799;
799: estado = 800;
800: estado = 801;
801: estado = 802;
802: estado = 803;
803: estado = 804;
804: estado = 805;
805: estado = 806;
806: estado = 807;
807: estado = 808;
808: estado = 809;
809: estado = 810;
810: estado = 811;
811: estado = 812;
812: estado = 813;
813: estado = 814;
814: estado = 815;
815: estado = 816;
816: estado = 817;
817: estado = 818;
818: estado = 819;
819: estado = 820;
820: estado = 821;
821: estado = 822;
822: estado = 823;
823: estado = 824;
824: estado = 825;
825: estado = 826;
826: estado = 827;
827: estado = 828;
828: estado = 829;
829: estado = 830;
830: estado = 831;
831: estado = 832;
832: estado = 833;
833: estado = 834;
834: estado = 835;
835: estado = 836;
836: estado = 837;
837: estado = 838;
838: estado = 839;
839: estado = 840;
840: estado = 841;
841: estado = 842;
842: estado = 843;
843: estado = 844;
844: estado = 845;
845: estado = 846;
846: estado = 847;
847: estado = 848;
848: estado = 849;
849: estado = 850;
850: estado = 851;
851: estado = 852;
852: estado = 853;
853: estado = 854;
854: estado = 855;
855: estado = 856;
856: estado = 857;
857: estado = 858;
858: estado = 859;
859: estado = 860;
860: estado = 861;
861: estado = 862;
862: estado = 863;
863: estado = 864;
864: estado = 865;
865: estado = 866;
866: estado = 867;
867: estado = 868;
868: estado = 869;
869: estado = 870;
870: estado = 871;
871: estado = 872;
872: estado = 873;
873: estado = 874;
874: estado = 875;
875: estado = 876;
876: estado = 877;
877: estado = 878;
878: estado = 879;
879: estado = 880;
880: estado = 881;
881: estado = 882;
882: estado = 883;
883: estado = 884;
884: estado = 885;
885: estado = 886;
886: estado = 887;
887: estado = 888;
888: estado = 889;
889: estado = 890;
890: estado = 891;
891: estado = 892;
892: estado = 893;
893: estado = 894;
894: estado = 895;
895: estado = 896;
896: estado = 897;
897: estado = 898;
898: estado = 899;
899: estado = 900;
900: estado = 901;
901: estado = 902;
902: estado = 903;
903: estado = 904;
904: estado = 905;
905: estado = 906;
906: estado = 907;
907: estado = 908;
908: estado = 909;
909: estado = 910;
910: estado = 911;
911: estado = 912;
912: estado = 913;
913: estado = 914;
914: estado = 915;
915: estado = 916;
916: estado = 917;
917: estado = 918;
918: estado = 919;
919: estado = 920;
920: estado = 921;
921: estado = 922;
922: estado = 923;
923: estado = 924;
924: estado = 925;
925: estado = 926;
926: estado = 927;
927: estado = 928;
928: estado = 929;
929: estado = 930;
930: estado = 931;
931: estado = 932;
932: estado = 933;
933: estado = 934;
934: estado = 935;
935: estado = 936;
936: estado = 937;
937: estado = 938;
938: estado = 939;
939: estado = 940;
940: estado = 941;
941: estado = 942;
942: estado = 943;
943: estado = 944;
944: estado = 945;
945: estado = 946;
946: estado = 947;
947: estado = 948;
948: estado = 949;
949: estado = 950;
950: estado = 951;
951: estado = 952;
952: estado = 953;
953: estado = 954;
954: estado = 955;
955: estado = 956;
956: estado = 957;
957: estado = 958;
958: estado = 959;
959: estado = 960;
960: estado = 961;
961: estado = 962;
962: estado = 963;
963: estado = 964;
964: estado = 965;
965: estado = 966;
966: estado = 967;
967: estado = 968;
968: estado = 969;
969: estado = 970;
970: estado = 971;
971: estado = 972;
972: estado = 973;
973: estado = 974;
974: estado = 975;
975: estado = 976;
976: estado = 977;
977: estado = 978;
978: estado = 979;
979: estado = 980;
980: estado = 981;
981: estado = 982;
982: estado = 983;
983: estado = 984;
984: estado = 985;
985: estado = 986;
986: estado = 987;
987: estado = 988;
988: estado = 989;
989: estado = 990;
990: estado = 991;
991: estado = 992;
992: estado = 993;
993: estado = 994;
994: estado = 995;
995: estado = 996;
996: estado = 997;
997: estado = 998;
998: estado = 999;
999: estado = 1000;
1000: estado = 1001;
1001: estado = 1002;
1002: estado = 1003;
1003: estado = 1004;
1004: estado = 1005;
1005: estado = 1006;
1006: estado = 1007;
1007: estado = 1008;
1008: estado = 1009;
1009: estado = 1010;
1010: estado = 1011;
1011: estado = 1012;
1012: estado = 1013;
1013: estado = 1014;
1014: estado = 1015;
1015: estado = 1016;
1016: estado = 1017;
1017: estado = 1018;
1018: estado = 1019;
1019: estado = 1020;
1020: estado = 1021;
1021: estado = 1022;
1022: estado = 1023;
1023: estado = 1024;
1024: estado = 1025;
1025: estado = 1026;
1026: estado = 1027;
1027: estado = 1028;
1028: estado = 1029;
1029: estado = 1030;
1030: estado = 1031;
1031: estado = 1032;
1032: estado = 1033;
1033: estado = 1034;
1034: estado = 1035;
1035: estado = 1036;
1036: estado = 1037;
1037: estado = 1038;
1038: estado = 1039;
1039: estado = 1040;
1040: estado = 1041;
1041: estado = 1042;
1042: estado = 1043;
1043: estado = 1044;
1044: estado = 1045;
1045: estado = 1046;
1046: estado = 1047;
1047: estado = 1048;
1048: estado = 1049;
1049: estado = 1050;
1050: estado = 1051;
1051: estado = 1052;
1052: estado = 1053;
1053: estado = 1054;
1054: estado = 1055;
1055: estado = 1056;
1056: estado = 1057;
1057: estado = 1058;
1058: estado = 1059;
1059: estado = 1060;
1060: estado = 1061;
1061: estado = 1062;
1062: estado = 1063;
1063: estado = 1064;
1064: estado = 1065;
1065: estado = 1066;
1066: estado = 1067;
1067: estado = 1068;
1068: estado = 1069;
1069: estado = 1070;
1070: estado = 1071;
1071: estado = 1072;
1072: estado = 1073;
1073: estado = 1074;
1074: estado = 1075;
1075: estado = 1076;
1076: estado = 1077;
1077: estado = 1078;
1078: estado = 1079;
1079: estado = 1080;
1080: estado = 1081;
1081: estado = 1082;
1082: estado = 1083;
1083: estado = 1084;
1084: estado = 1085;
1085: estado = 1086;
1086: estado = 1087;
1087: estado = 1088;
1088: estado = 1089;
1089: estado = 1090;
1090: estado = 1091;
1091: estado = 1092;
1092: estado = 1093;
1093: estado = 1094;
1094: estado = 1095;
1095: estado = 1096;
1096: estado = 1097;
1097: estado = 1098;
1098: estado = 1099;
1099: estado = 1100;
1100: estado = 1101;
1101: estado = 1102;
1102: estado = 1103;
1103: estado = 1104;
1104: estado = 1105;
1105: estado = 1106;
1106: estado = 1107;
1107: estado = 1108;
1108: estado = 1109;
1109: estado = 1110;
1110: estado = 1111;
1111: estado = 1112;
1112: estado = 1113;
1113: estado = 1114;
1114: estado = 1115;
1115: estado = 1116;
1116: estado = 1117;
1117: estado = 1118;
1118: estado = 1119;
1119: estado = 1120;
1120: estado = 1121;
1121: estado = 1122;
1122: estado = 1123;
1123: estado = 1124;
1124: estado = 1125;
1125: estado = 1126;
1126: estado = 1127;
1127: estado = 1128;
1128: estado = 1129;
1129: estado = 1130;
1130: estado = 1131;
1131: estado = 1132;
1132: estado = 1133;
1133: estado = 1134;
1134: estado = 1135;
1135: estado = 1136;
1136: estado = 1137;
1137: estado = 1138;
1138: estado = 1139;
1139: estado = 1140;
1140: estado = 1141;
1141: estado = 1142;
1142: estado = 1143;
1143: estado = 1144;
1144: estado = 1145;
1145: estado = 1146;
1146: estado = 1147;
1147: estado = 1148;
1148: estado = 1149;
1149: estado = 1150;
1150: estado = 1151;
1151: estado = 1152;
1152: estado = 1153;
1153: estado = 1154;
1154: estado = 1155;
1155: estado = 1156;
1156: estado = 1157;
1157: estado = 1158;
1158: estado = 1159;
1159: estado = 1160;
1160: estado = 1161;
1161: estado = 1162;
1162: estado = 1163;
1163: estado = 1164;
1164: estado = 1165;
1165: estado = 1166;
1166: estado = 1167;
1167: estado = 1168;
1168: estado = 1169;
1169: estado = 1170;
1170: estado = 1171;
1171: estado = 1172;
1172: estado = 1173;
1173: estado = 1174;
1174: estado = 1175;
1175: estado = 1176;
1176: estado = 1177;
1177: estado = 1178;
1178: estado = 1179;
1179: estado = 1180;
1180: estado = 1181;
1181: estado = 1182;
1182: estado = 1183;
1183: estado = 1184;
1184: estado = 1185;
1185: estado = 1186;
1186: estado = 1187;
1187: estado = 1188;
1188: estado = 1189;
1189: estado = 1190;
1190: estado = 1191;
1191: estado = 1192;
1192: estado = 1193;
1193: estado = 1194;
1194: estado = 1195;
1195: estado = 1196;
1196: estado = 1197;
1197: estado = 1198;
1198: estado = 1199;
1199: estado = 1200;
1200: estado = 1201;
1201: estado = 1202;
1202: estado = 1203;
1203: estado = 1204;
1204: estado = 1205;
1205: estado = 1206;
1206: estado = 1207;
1207: estado = 1208;
1208: estado = 1209;
1209: estado = 1210;
1210: estado = 1211;
1211: estado = 1212;
1212: estado = 1213;
1213: estado = 1214;
1214: estado = 1215;
1215: estado = 1216;
1216: estado = 1217;
1217: estado = 1218;
1218: estado = 1219;
1219: estado = 1220;
1220: estado = 1221;
1221: estado = 1222;
1222: estado = 1223;
1223: estado = 1224;
1224: estado = 1225;
1225: estado = 1226;
1226: estado = 1227;
1227: estado = 1228;
1228: estado = 1229;
1229: estado = 1230;
1230: estado = 1231;
1231: estado = 1232;
1232: estado = 1233;
1233: estado = 1234;
1234: estado = 1235;
1235: estado = 1236;
1236: estado = 1237;
1237: estado = 1238;
1238: estado = 1239;
1239: estado = 1240;
1240: estado = 1241;
1241: estado = 1242;
1242: estado = 1243;
1243: estado = 1244;
1244: estado = 1245;
1245: estado = 1246;
1246: estado = 1247;
1247: estado = 1248;
1248: estado = 1249;
1249: estado = 1250;
1250: estado = 1251;
1251: estado = 1252;
1252: estado = 1253;
1253: estado = 1254;
1254: estado = 1255;
1255: estado = 1256;
1256: estado = 1257;
1257: estado = 1258;
1258: estado = 1259;
1259: estado = 1260;
1260: estado = 1261;
1261: estado = 1262;
1262: estado = 1263;
1263: estado = 1264;
1264: estado = 1265;
1265: estado = 1266;
1266: estado = 1267;
1267: estado = 1268;
1268: estado = 1269;
1269: estado = 1270;
1270: estado = 1271;
1271: estado = 1272;
1272: estado = 1273;
1273: estado = 1274;
1274: estado = 1275;
1275: estado = 1276;
1276: estado = 1277;
1277: estado = 1278;
1278: estado = 1279;
1279: estado = 1280;
1280: estado = 1281;
1281: estado = 1282;
1282: estado = 1283;
1283: estado = 1284;
1284: estado = 1285;
1285: estado = 1286;
1286: estado = 1287;
1287: estado = 1288;
1288: estado = 1289;
1289: estado = 1290;
1290: estado = 1291;
1291: estado = 1292;
1292: estado = 1293;
1293: estado = 1294;
1294: estado = 1295;
1295: estado = 1296;
1296: estado = 1297;
1297: estado = 1298;
1298: estado = 1299;
1299: estado = 1300;
1300: estado = 1301;
1301: estado = 1302;
1302: estado = 1303;
1303: estado = 1304;
1304: estado = 1305;
1305: estado = 1306;
1306: estado = 1307;
1307: estado = 1308;
1308: estado = 1309;
1309: estado = 1310;
1310: estado = 1311;
1311: estado = 1312;
1312: estado = 1313;
1313: estado = 1314;
1314: estado = 1315;
1315: estado = 1316;
1316: estado = 1317;
1317: estado = 1318;
1318: estado = 1319;
1319: estado = 1320;
1320: estado = 1321;
1321: estado = 1322;
1322: estado = 1323;
1323: estado = 1324;
1324: estado = 1325;
1325: estado = 1326;
1326: estado = 1327;
1327: estado = 1328;
1328: estado = 1329;
1329: estado = 1330;
1330: estado = 1331;
1331: estado = 1332;
1332: estado = 1333;
1333: estado = 1334;
1334: estado = 1335;
1335: estado = 1336;
1336: estado = 1337;
1337: estado = 1338;
1338: estado = 1339;
1339: estado = 1340;
1340: estado = 1341;
1341: estado = 1342;
1342: estado = 1343;
1343: estado = 1344;
1344: estado = 1345;
1345: estado = 1346;
1346: estado = 1347;
1347: estado = 1348;
1348: estado = 1349;
1349: estado = 1350;
1350: estado = 1351;
1351: estado = 1352;
1352: estado = 1353;
1353: estado = 1354;
1354: estado = 1355;
1355: estado = 1356;
1356: estado = 1357;
1357: estado = 1358;
1358: estado = 1359;
1359: estado = 1360;
1360: estado = 1361;
1361: estado = 1362;
1362: estado = 1363;
1363: estado = 1364;
1364: estado = 1365;
1365: estado = 1366;
1366: estado = 1367;
1367: estado = 1368;
1368: estado = 1369;
1369: estado = 1370;
1370: estado = 1371;
1371: estado = 1372;
1372: estado = 1373;
1373: estado = 1374;
1374: estado = 1375;
1375: estado = 1376;
1376: estado = 1377;
1377: estado = 1378;
1378: estado = 1379;
1379: estado = 1380;
1380: estado = 1381;
1381: estado = 1382;
1382: estado = 1383;
1383: estado = 1384;
1384: estado = 1385;
1385: estado = 1386;
1386: estado = 1387;
1387: estado = 1388;
1388: estado = 1389;
1389: estado = 1390;
1390: estado = 1391;
1391: estado = 1392;
1392: estado = 1393;
1393: estado = 1394;
1394: estado = 1395;
1395: estado = 1396;
1396: estado = 1397;
1397: estado = 1398;
1398: estado = 1399;
1399: estado = 1400;
1400: estado = 1401;
1401: estado = 1402;
1402: estado = 1403;
1403: estado = 1404;
1404: estado = 1405;
1405: estado = 1406;
1406: estado = 1407;
1407: estado = 1408;
1408: estado = 1409;
1409: estado = 1410;
1410: estado = 1411;
1411: estado = 1412;
1412: estado = 1413;
1413: estado = 1414;
1414: estado = 1415;
1415: estado = 1416;
1416: estado = 1417;
1417: estado = 1418;
1418: estado = 1419;
1419: estado = 1420;
1420: estado = 1421;
1421: estado = 1422;
1422: estado = 1423;
1423: estado = 1424;
1424: estado = 1425;
1425: estado = 1426;
1426: estado = 1427;
1427: estado = 1428;
1428: estado = 1429;
1429: estado = 1430;
1430: estado = 1431;
1431: estado = 1432;
1432: estado = 1433;
1433: estado = 1434;
1434: estado = 1435;
1435: estado = 1436;
1436: estado = 1437;
1437: estado = 1438;
1438: estado = 1439;
1439: estado = 1440;
1440: estado = 1441;
1441: estado = 1442;
1442: estado = 1443;
1443: estado = 1444;
1444: estado = 1445;
1445: estado = 1446;
1446: estado = 1447;
1447: estado = 1448;
1448: estado = 1449;
1449: estado = 1450;
1450: estado = 1451;
1451: estado = 1452;
1452: estado = 1453;
1453: estado = 1454;
1454: estado = 1455;
1455: estado = 1456;
1456: estado = 1457;
1457: estado = 1458;
1458: estado = 1459;
1459: estado = 1460;
1460: estado = 1461;
1461: estado = 1462;
1462: estado = 1463;
1463: estado = 1464;
1464: estado = 1465;
1465: estado = 1466;
1466: estado = 1467;
1467: estado = 1468;
1468: estado = 1469;
1469: estado = 1470;
1470: estado = 1471;
1471: estado = 1472;
1472: estado = 1473;
1473: estado = 1474;
1474: estado = 1475;
1475: estado = 1476;
1476: estado = 1477;
1477: estado = 1478;
1478: estado = 1479;
1479: estado = 1480;
1480: estado = 1481;
1481: estado = 1482;
1482: estado = 1483;
1483: estado = 1484;
1484: estado = 1485;
1485: estado = 1486;
1486: estado = 1487;
1487: estado = 1488;
1488: estado = 1489;
1489: estado = 1490;
1490: estado = 1491;
1491: estado = 1492;
1492: estado = 1493;
1493: estado = 1494;
1494: estado = 1495;
1495: estado = 1496;
1496: estado = 1497;
1497: estado = 1498;
1498: estado = 1499;
1499: estado = 1500;
1500: estado = 1501;
1501: estado = 1502;
1502: estado = 1503;
1503: estado = 1504;
1504: estado = 1505;
1505: estado = 1506;
1506: estado = 1507;
1507: estado = 1508;
1508: estado = 1509;
1509: estado = 1510;
1510: estado = 1511;
1511: estado = 1512;
1512: estado = 1513;
1513: estado = 1514;
1514: estado = 1515;
1515: estado = 1516;
1516: estado = 1517;
1517: estado = 1518;
1518: estado = 1519;
1519: estado = 1520;
1520: estado = 1521;
1521: estado = 1522;
1522: estado = 1523;
1523: estado = 1524;
1524: estado = 1525;
1525: estado = 1526;
1526: estado = 1527;
1527: estado = 1528;
1528: estado = 1529;
1529: estado = 1530;
1530: estado = 1531;
1531: estado = 1532;
1532: estado = 1533;
1533: estado = 1534;
1534: estado = 1535;
1535: estado = 1536;
1536: estado = 1537;
1537: estado = 1538;
1538: estado = 1539;
1539: estado = 1540;
1540: estado = 1541;
1541: estado = 1542;
1542: estado = 1543;
1543: estado = 1544;
1544: estado = 1545;
1545: estado = 1546;
1546: estado = 1547;
1547: estado = 1548;
1548: estado = 1549;
1549: estado = 1550;
1550: estado = 1551;
1551: estado = 1552;
1552: estado = 1553;
1553: estado = 1554;
1554: estado = 1555;
1555: estado = 1556;
1556: estado = 1557;
1557: estado = 1558;
1558: estado = 1559;
1559: estado = 1560;
1560: estado = 1561;
1561: estado = 1562;
1562: estado = 1563;
1563: estado = 1564;
1564: estado = 1565;
1565: estado = 1566;
1566: estado = 1567;
1567: estado = 1568;
1568: estado = 1569;
1569: estado = 1570;
1570: estado = 1571;
1571: estado = 1572;
1572: estado = 1573;
1573: estado = 1574;
1574: estado = 1575;
1575: estado = 1576;
1576: estado = 1577;
1577: estado = 1578;
1578: estado = 1579;
1579: estado = 1580;
1580: estado = 1581;
1581: estado = 1582;
1582: estado = 1583;
1583: estado = 1584;
1584: estado = 1585;
1585: estado = 1586;
1586: estado = 1587;
1587: estado = 1588;
1588: estado = 1589;
1589: estado = 1590;
1590: estado = 1591;
1591: estado = 1592;
1592: estado = 1593;
1593: estado = 1594;
1594: estado = 1595;
1595: estado = 1596;
1596: estado = 1597;
1597: estado = 1598;
1598: estado = 1599;
1599: estado = 1600;
1600: estado = 1601;
1601: estado = 1602;
1602: estado = 1603;
1603: estado = 1604;
1604: estado = 1605;
1605: estado = 1606;
1606: estado = 1607;
1607: estado = 1608;
1608: estado = 1609;
1609: estado = 1610;
1610: estado = 1611;
1611: estado = 1612;
1612: estado = 1613;
1613: estado = 1614;
1614: estado = 1615;
1615: estado = 1616;
1616: estado = 1617;
1617: estado = 1618;
1618: estado = 1619;
1619: estado = 1620;
1620: estado = 1621;
1621: estado = 1622;
1622: estado = 1623;
1623: estado = 1624;
1624: estado = 1625;
1625: estado = 1626;
1626: estado = 1627;
1627: estado = 1628;
1628: estado = 1629;
1629: estado = 1630;
1630: estado = 1631;
1631: estado = 1632;
1632: estado = 1633;
1633: estado = 1634;
1634: estado = 1635;
1635: estado = 1636;
1636: estado = 1637;
1637: estado = 1638;
1638: estado = 1639;
1639: estado = 1640;
1640: estado = 1641;
1641: estado = 1642;
1642: estado = 1643;
1643: estado = 1644;
1644: estado = 1645;
1645: estado = 1646;
1646: estado = 1647;
1647: estado = 1648;
1648: estado = 1649;
1649: estado = 1650;
1650: estado = 1651;
1651: estado = 1652;
1652: estado = 1653;
1653: estado = 1654;
1654: estado = 1655;
1655: estado = 1656;
1656: estado = 1657;
1657: estado = 1658;
1658: estado = 1659;
1659: estado = 1660;
1660: estado = 1661;
1661: estado = 1662;
1662: estado = 1663;
1663: estado = 1664;
1664: estado = 1665;
1665: estado = 1666;
1666: estado = 1667;
1667: estado = 1668;
1668: estado = 1669;
1669: estado = 1670;
1670: estado = 1671;
1671: estado = 1672;
1672: estado = 1673;
1673: estado = 1674;
1674: estado = 1675;
1675: estado = 1676;
1676: estado = 1677;
1677: estado = 1678;
1678: estado = 1679;
1679: estado = 1680;
1680: estado = 1681;
1681: estado = 1682;
1682: estado = 1683;
1683: estado = 1684;
1684: estado = 1685;
1685: estado = 1686;
1686: estado = 1687;
1687: estado = 1688;
1688: estado = 1689;
1689: estado = 1690;
1690: estado = 1691;
1691: estado = 1692;
1692: estado = 1693;
1693: estado = 1694;
1694: estado = 1695;
1695: estado = 1696;
1696: estado = 1697;
1697: estado = 1698;
1698: estado = 1699;
1699: estado = 1700;
1700: estado = 1701;
1701: estado = 1702;
1702: estado = 1703;
1703: estado = 1704;
1704: estado = 1705;
1705: estado = 1706;
1706: estado = 1707;
1707: estado = 1708;
1708: estado = 1709;
1709: estado = 1710;
1710: estado = 1711;
1711: estado = 1712;
1712: estado = 1713;
1713: estado = 1714;
1714: estado = 1715;
1715: estado = 1716;
1716: estado = 1717;
1717: estado = 1718;
1718: estado = 1719;
1719: estado = 1720;
1720: estado = 1721;
1721: estado = 1722;
1722: estado = 1723;
1723: estado = 1724;
1724: estado = 1725;
1725: estado = 1726;
1726: estado = 1727;
1727: estado = 1728;
1728: estado = 1729;
1729: estado = 1730;
1730: estado = 1731;
1731: estado = 1732;
1732: estado = 1733;
1733: estado = 1734;
1734: estado = 1735;
1735: estado = 1736;
1736: estado = 1737;
1737: estado = 1738;
1738: estado = 1739;
1739: estado = 1740;
1740: estado = 1741;
1741: estado = 1742;
1742: estado = 1743;
1743: estado = 1744;
1744: estado = 1745;
1745: estado = 1746;
1746: estado = 1747;
1747: estado = 1748;
1748: estado = 1749;
1749: estado = 1750;
1750: estado = 1751;
1751: estado = 1752;
1752: estado = 1753;
1753: estado = 1754;
1754: estado = 1755;
1755: estado = 1756;
1756: estado = 1757;
1757: estado = 1758;
1758: estado = 1759;
1759: estado = 1760;
1760: estado = 1761;
1761: estado = 1762;
1762: estado = 1763;
1763: estado = 1764;
1764: estado = 1765;
1765: estado = 1766;
1766: estado = 1767;
1767: estado = 1768;
1768: estado = 1769;
1769: estado = 1770;
1770: estado = 1771;
1771: estado = 1772;
1772: estado = 1773;
1773: estado = 1774;
1774: estado = 1775;
1775: estado = 1776;
1776: estado = 1777;
1777: estado = 1778;
1778: estado = 1779;
1779: estado = 1780;
1780: estado = 1781;
1781: estado = 1782;
1782: estado = 1783;
1783: estado = 1784;
1784: estado = 1785;
1785: estado = 1786;
1786: estado = 1787;
1787: estado = 1788;
1788: estado = 1789;
1789: estado = 1790;
1790: estado = 1791;
1791: estado = 1792;
1792: estado = 1793;
1793: estado = 1794;
1794: estado = 1795;
1795: estado = 1796;
1796: estado = 1797;
1797: estado = 1798;
1798: estado = 1799;
1799: estado = 1800;
1800: estado = 1801;
1801: estado = 1802;
1802: estado = 1803;
1803: estado = 1804;
1804: estado = 1805;
1805: estado = 1806;
1806: estado = 1807;
1807: estado = 1808;
1808: estado = 1809;
1809: estado = 1810;
1810: estado = 1811;
1811: estado = 1812;
1812: estado = 1813;
1813: estado = 1814;
1814: estado = 1815;
1815: estado = 1816;
1816: estado = 1817;
1817: estado = 1818;
1818: estado = 1819;
1819: estado = 1820;
1820: estado = 1821;
1821: estado = 1822;
1822: estado = 1823;
1823: estado = 1824;
1824: estado = 1825;
1825: estado = 1826;
1826: estado = 1827;
1827: estado = 1828;
1828: estado = 1829;
1829: estado = 1830;
1830: estado = 1831;
1831: estado = 1832;
1832: estado = 1833;
1833: estado = 1834;
1834: estado = 1835;
1835: estado = 1836;
1836: estado = 1837;
1837: estado = 1838;
1838: estado = 1839;
1839: estado = 1840;
1840: estado = 1841;
1841: estado = 1842;
1842: estado = 1843;
1843: estado = 1844;
1844: estado = 1845;
1845: estado = 1846;
1846: estado = 1847;
1847: estado = 1848;
1848: estado = 1849;
1849: estado = 1850;
1850: estado = 1851;
1851: estado = 1852;
1852: estado = 1853;
1853: estado = 1854;
1854: estado = 1855;
1855: estado = 1856;
1856: estado = 1857;
1857: estado = 1858;
1858: estado = 1859;
1859: estado = 1860;
1860: estado = 1861;
1861: estado = 1862;
1862: estado = 1863;
1863: estado = 1864;
1864: estado = 1865;
1865: estado = 1866;
1866: estado = 1867;
1867: estado = 1868;
1868: estado = 1869;
1869: estado = 1870;
1870: estado = 1871;
1871: estado = 1872;
1872: estado = 1873;
1873: estado = 1874;
1874: estado = 1875;
1875: estado = 1876;
1876: estado = 1877;
1877: estado = 1878;
1878: estado = 1879;
1879: estado = 1880;
1880: estado = 1881;
1881: estado = 1882;
1882: estado = 1883;
1883: estado = 1884;
1884: estado = 1885;
1885: estado = 1886;
1886: estado = 1887;
1887: estado = 1888;
1888: estado = 1889;
1889: estado = 1890;
1890: estado = 1891;
1891: estado = 1892;
1892: estado = 1893;
1893: estado = 1894;
1894: estado = 1895;
1895: estado = 1896;
1896: estado = 1897;
1897: estado = 1898;
1898: estado = 1899;
1899: estado = 1900;
1900: estado = 1901;
1901: estado = 1902;
1902: estado = 1903;
1903: estado = 1904;
1904: estado = 1905;
1905: estado = 1906;
1906: estado = 1907;
1907: estado = 1908;
1908: estado = 1909;
1909: estado = 1910;
1910: estado = 1911;
1911: estado = 1912;
1912: estado = 1913;
1913: estado = 1914;
1914: estado = 1915;
1915: estado = 1916;
1916: estado = 1917;
1917: estado = 1918;
1918: estado = 1919;
1919: estado = 1920;
1920: estado = 1921;
1921: estado = 1922;
1922: estado = 1923;
1923: estado = 1924;
1924: estado = 1925;
1925: estado = 1926;
1926: estado = 1927;
1927: estado = 1928;
1928: estado = 1929;
1929: estado = 1930;
1930: estado = 1931;
1931: estado = 1932;
1932: estado = 1933;
1933: estado = 1934;
1934: estado = 1935;
1935: estado = 1936;
1936: estado = 1937;
1937: estado = 1938;
1938: estado = 1939;
1939: estado = 1940;
1940: estado = 1941;
1941: estado = 1942;
1942: estado = 1943;
1943: estado = 1944;
1944: estado = 1945;
1945: estado = 1946;
1946: estado = 1947;
1947: estado = 1948;
1948: estado = 1949;
1949: estado = 1950;
1950: estado = 1951;
1951: estado = 1952;
1952: estado = 1953;
1953: estado = 1954;
1954: estado = 1955;
1955: estado = 1956;
1956: estado = 1957;
1957: estado = 1958;
1958: estado = 1959;
1959: estado = 1960;
1960: estado = 1961;
1961: estado = 1962;
1962: estado = 1963;
1963: estado = 1964;
1964: estado = 1965;
1965: estado = 1966;
1966: estado = 1967;
1967: estado = 1968;
1968: estado = 1969;
1969: estado = 1970;
1970: estado = 1971;
1971: estado = 1972;
1972: estado = 1973;
1973: estado = 1974;
1974: estado = 1975;
1975: estado = 1976;
1976: estado = 1977;
1977: estado = 1978;
1978: estado = 1979;
1979: estado = 1980;
1980: estado = 1981;
1981: estado = 1982;
1982: estado = 1983;
1983: estado = 1984;
1984: estado = 1985;
1985: estado = 1986;
1986: estado = 1987;
1987: estado = 1988;
1988: estado = 1989;
1989: estado = 1990;
1990: estado = 1991;
1991: estado = 1992;
1992: estado = 1993;
1993: estado = 1994;
1994: estado = 1995;
1995: estado = 1996;
1996: estado = 1997;
1997: estado = 1998;
1998: estado = 1999;
1999: estado = 2000;
2000: estado = 2001;
2001: estado = 2002;
2002: estado = 2003;
2003: estado = 2004;
2004: estado = 2005;
2005: estado = 2006;
2006: estado = 2007;
2007: estado = 2008;
2008: estado = 2009;
2009: estado = 2010;
2010: estado = 2011;
2011: estado = 2012;
2012: estado = 2013;
2013: estado = 2014;
2014: estado = 2015;
2015: estado = 2016;
2016: estado = 2017;
2017: estado = 2018;
2018: estado = 2019;
2019: estado = 2020;
2020: estado = 2021;
2021: estado = 2022;
2022: estado = 2023;
2023: estado = 2024;
2024: estado = 2025;
2025: estado = 2026;
2026: estado = 2027;
2027: estado = 2028;
2028: estado = 2029;
2029: estado = 2030;
2030: estado = 2031;
2031: estado = 2032;
2032: estado = 2033;
2033: estado = 2034;
2034: estado = 2035;
2035: estado = 2036;
2036: estado = 2037;
2037: estado = 2038;
2038: estado = 2039;
2039: estado = 2040;
2040: estado = 2041;
2041: estado = 2042;
2042: estado = 2043;
2043: estado = 2044;
2044: estado = 2045;
2045: estado = 2046;
2046: estado = 2047;
2047: estado = 2048;
2048: estado = 2049;
2049: estado = 2050;
2050: estado = 2051;
2051: estado = 2052;
2052: estado = 2053;
2053: estado = 2054;
2054: estado = 2055;
2055: estado = 2056;
2056: estado = 2057;
2057: estado = 2058;
2058: estado = 2059;
2059: estado = 2060;
2060: estado = 2061;
2061: estado = 2062;
2062: estado = 2063;
2063: estado = 2064;
2064: estado = 2065;
2065: estado = 2066;
2066: estado = 2067;
2067: estado = 2068;
2068: estado = 2069;
2069: estado = 2070;
2070: estado = 2071;
2071: estado = 2072;
2072: estado = 2073;
2073: estado = 2074;
2074: estado = 2075;
2075: estado = 2076;
2076: estado = 2077;
2077: estado = 2078;
2078: estado = 2079;
2079: estado = 2080;
2080: estado = 2081;
2081: estado = 2082;
2082: estado = 2083;
2083: estado = 2084;
2084: estado = 2085;
2085: estado = 2086;
2086: estado = 2087;
2087: estado = 2088;
2088: estado = 2089;
2089: estado = 2090;
2090: estado = 2091;
2091: estado = 2092;
2092: estado = 2093;
2093: estado = 2094;
2094: estado = 2095;
2095: estado = 2096;
2096: estado = 2097;
2097: estado = 2098;
2098: estado = 2099;
2099: estado = 2100;
2100: estado = 2101;
2101: estado = 2102;
2102: estado = 2103;
2103: estado = 2104;
2104: estado = 2105;
2105: estado = 2106;
2106: estado = 2107;
2107: estado = 2108;
2108: estado = 2109;
2109: estado = 2110;
2110: estado = 2111;
2111: estado = 2112;
2112: estado = 2113;
2113: estado = 2114;
2114: estado = 2115;
2115: estado = 2116;
2116: estado = 2117;
2117: estado = 2118;
2118: estado = 2119;
2119: estado = 2120;
2120: estado = 2121;
2121: estado = 2122;
2122: estado = 2123;
2123: estado = 2124;
2124: estado = 2125;
2125: estado = 2126;
2126: estado = 2127;
2127: estado = 2128;
2128: estado = 2129;
2129: estado = 2130;
2130: estado = 2131;
2131: estado = 2132;
2132: estado = 2133;
2133: estado = 2134;
2134: estado = 2135;
2135: estado = 2136;
2136: estado = 2137;
2137: estado = 2138;
2138: estado = 2139;
2139: estado = 2140;
2140: estado = 2141;
2141: estado = 2142;
2142: estado = 2143;
2143: estado = 2144;
2144: estado = 2145;
2145: estado = 2146;
2146: estado = 2147;
2147: estado = 2148;
2148: estado = 2149;
2149: estado = 2150;
2150: estado = 2151;
2151: estado = 2152;
2152: estado = 2153;
2153: estado = 2154;
2154: estado = 2155;
2155: estado = 2156;
2156: estado = 2157;
2157: estado = 2158;
2158: estado = 2159;
2159: estado = 2160;
2160: estado = 2161;
2161: estado = 2162;
2162: estado = 2163;
2163: estado = 2164;
2164: estado = 2165;
2165: estado = 2166;
2166: estado = 2167;
2167: estado = 2168;
2168: estado = 2169;
2169: estado = 2170;
2170: estado = 2171;
2171: estado = 2172;
2172: estado = 2173;
2173: estado = 2174;
2174: estado = 2175;
2175: estado = 2176;
2176: estado = 2177;
2177: estado = 2178;
2178: estado = 2179;
2179: estado = 2180;
2180: estado = 2181;
2181: estado = 2182;
2182: estado = 2183;
2183: estado = 2184;
2184: estado = 2185;
2185: estado = 2186;
2186: estado = 2187;
2187: estado = 2188;
2188: estado = 2189;
2189: estado = 2190;
2190: estado = 2191;
2191: estado = 2192;
2192: estado = 2193;
2193: estado = 2194;
2194: estado = 2195;
2195: estado = 2196;
2196: estado = 2197;
2197: estado = 2198;
2198: estado = 2199;
2199: estado = 2200;
2200: estado = 2201;
2201: estado = 2202;
2202: estado = 2203;
2203: estado = 2204;
2204: estado = 2205;
2205: estado = 2206;
2206: estado = 2207;
2207: estado = 2208;
2208: estado = 2209;
2209: estado = 2210;
2210: estado = 2211;
2211: estado = 2212;
2212: estado = 2213;
2213: estado = 2214;
2214: estado = 2215;
2215: estado = 2216;
2216: estado = 2217;
2217: estado = 2218;
2218: estado = 2219;
2219: estado = 2220;
2220: estado = 2221;
2221: estado = 2222;
2222: estado = 2223;
2223: estado = 2224;
2224: estado = 2225;
2225: estado = 2226;
2226: estado = 2227;
2227: estado = 2228;
2228: estado = 2229;
2229: estado = 2230;
2230: estado = 2231;
2231: estado = 2232;
2232: estado = 2233;
2233: estado = 2234;
2234: estado = 2235;
2235: estado = 2236;
2236: estado = 2237;
2237: estado = 2238;
2238: estado = 2239;
2239: estado = 2240;
2240: estado = 2241;
2241: estado = 2242;
2242: estado = 2243;
2243: estado = 2244;
2244: estado = 2245;
2245: estado = 2246;
2246: estado = 2247;
2247: estado = 2248;
2248: estado = 2249;
2249: estado = 2250;
2250: estado = 2251;
2251: estado = 2252;
2252: estado = 2253;
2253: estado = 2254;
2254: estado = 2255;
2255: estado = 2256;
2256: estado = 2257;
2257: estado = 2258;
2258: estado = 2259;
2259: estado = 2260;
2260: estado = 2261;
2261: estado = 2262;
2262: estado = 2263;
2263: estado = 2264;
2264: estado = 2265;
2265: estado = 2266;
2266: estado = 2267;
2267: estado = 2268;
2268: estado = 2269;
2269: estado = 2270;
2270: estado = 2271;
2271: estado = 2272;
2272: estado = 2273;
2273: estado = 2274;
2274: estado = 2275;
2275: estado = 2276;
2276: estado = 2277;
2277: estado = 2278;
2278: estado = 2279;
2279: estado = 2280;
2280: estado = 2281;
2281: estado = 2282;
2282: estado = 2283;
2283: estado = 2284;
2284: estado = 2285;
2285: estado = 2286;
2286: estado = 2287;
2287: estado = 2288;
2288: estado = 2289;
2289: estado = 2290;
2290: estado = 2291;
2291: estado = 2292;
2292: estado = 2293;
2293: estado = 2294;
2294: estado = 2295;
2295: estado = 2296;
2296: estado = 2297;
2297: estado = 2298;
2298: estado = 2299;
2299: estado = 2300;
2300: estado = 2301;
2301: estado = 2302;
2302: estado = 2303;
2303: estado = 2304;
2304: estado = 2305;
2305: estado = 2306;
2306: estado = 2307;
2307: estado = 2308;
2308: estado = 2309;
2309: estado = 2310;
2310: estado = 2311;
2311: estado = 2312;
2312: estado = 2313;
2313: estado = 2314;
2314: estado = 2315;
2315: estado = 2316;
2316: estado = 2317;
2317: estado = 2318;
2318: estado = 2319;
2319: estado = 2320;
2320: estado = 2321;
2321: estado = 2322;
2322: estado = 2323;
2323: estado = 2324;
2324: estado = 2325;
2325: estado = 2326;
2326: estado = 2327;
2327: estado = 2328;
2328: estado = 2329;
2329: estado = 2330;
2330: estado = 2331;
2331: estado = 2332;
2332: estado = 2333;
2333: estado = 2334;
2334: estado = 2335;
2335: estado = 2336;
2336: estado = 2337;
2337: estado = 2338;
2338: estado = 2339;
2339: estado = 2340;
2340: estado = 2341;
2341: estado = 2342;
2342: estado = 2343;
2343: estado = 2344;
2344: estado = 2345;
2345: estado = 2346;
2346: estado = 2347;
2347: estado = 2348;
2348: estado = 2349;
2349: estado = 2350;
2350: estado = 2351;
2351: estado = 2352;
2352: estado = 2353;
2353: estado = 2354;
2354: estado = 2355;
2355: estado = 2356;
2356: estado = 2357;
2357: estado = 2358;
2358: estado = 2359;
2359: estado = 2360;
2360: estado = 2361;
2361: estado = 2362;
2362: estado = 2363;
2363: estado = 2364;
2364: estado = 2365;
2365: estado = 2366;
2366: estado = 2367;
2367: estado = 2368;
2368: estado = 2369;
2369: estado = 2370;
2370: estado = 2371;
2371: estado = 2372;
2372: estado = 2373;
2373: estado = 2374;
2374: estado = 2375;
2375: estado = 2376;
2376: estado = 2377;
2377: estado = 2378;
2378: estado = 2379;
2379: estado = 2380;
2380: estado = 2381;
2381: estado = 2382;
2382: estado = 2383;
2383: estado = 2384;
2384: estado = 2385;
2385: estado = 2386;
2386: estado = 2387;
2387: estado = 2388;
2388: estado = 2389;
2389: estado = 2390;
2390: estado = 2391;
2391: estado = 2392;
2392: estado = 2393;
2393: estado = 2394;
2394: estado = 2395;
2395: estado = 2396;
2396: estado = 2397;
2397: estado = 2398;
2398: estado = 2399;
2399: estado = 2400;
2400: estado = 2401;
2401: estado = 2402;
2402: estado = 2403;
2403: estado = 2404;
2404: estado = 2405;
2405: estado = 2406;
2406: estado = 2407;
2407: estado = 2408;
2408: estado = 2409;
2409: estado = 2410;
2410: estado = 2411;
2411: estado = 2412;
2412: estado = 2413;
2413: estado = 2414;
2414: estado = 2415;
2415: estado = 2416;
2416: estado = 2417;
2417: estado = 2418;
2418: estado = 2419;
2419: estado = 2420;
2420: estado = 2421;
2421: estado = 2422;
2422: estado = 2423;
2423: estado = 2424;
2424: estado = 2425;
2425: estado = 2426;
2426: estado = 2427;
2427: estado = 2428;
2428: estado = 2429;
2429: estado = 2430;
2430: estado = 2431;
2431: estado = 2432;
2432: estado = 2433;
2433: estado = 2434;
2434: estado = 2435;
2435: estado = 2436;
2436: estado = 2437;
2437: estado = 2438;
2438: estado = 2439;
2439: estado = 2440;
2440: estado = 2441;
2441: estado = 2442;
2442: estado = 2443;
2443: estado = 2444;
2444: estado = 2445;
2445: estado = 2446;
2446: estado = 2447;
2447: estado = 2448;
2448: estado = 2449;
2449: estado = 2450;
2450: estado = 2451;
2451: estado = 2452;
2452: estado = 2453;
2453: estado = 2454;
2454: estado = 2455;
2455: estado = 2456;
2456: estado = 2457;
2457: estado = 2458;
2458: estado = 2459;
2459: estado = 2460;
2460: estado = 2461;
2461: estado = 2462;
2462: estado = 2463;
2463: estado = 2464;
2464: estado = 2465;
2465: estado = 2466;
2466: estado = 2467;
2467: estado = 2468;
2468: estado = 2469;
2469: estado = 2470;
2470: estado = 2471;
2471: estado = 2472;
2472: estado = 2473;
2473: estado = 2474;
2474: estado = 2475;
2475: estado = 2476;
2476: estado = 2477;
2477: estado = 2478;
2478: estado = 2479;
2479: estado = 2480;
2480: estado = 2481;
2481: estado = 2482;
2482: estado = 2483;
2483: estado = 2484;
2484: estado = 2485;
2485: estado = 2486;
2486: estado = 2487;
2487: estado = 2488;
2488: estado = 2489;
2489: estado = 2490;
2490: estado = 2491;
2491: estado = 2492;
2492: estado = 2493;
2493: estado = 2494;
2494: estado = 2495;
2495: estado = 2496;
2496: estado = 2497;
2497: estado = 2498;
2498: estado = 2499;
2499: estado = 2500;
2500: estado = 2501;
2501: estado = 2502;
2502: estado = 2503;
2503: estado = 2504;
2504: estado = 2505;
2505: estado = 2506;
2506: estado = 2507;
2507: estado = 2508;
2508: estado = 2509;
2509: estado = 2510;
2510: estado = 2511;
2511: estado = 2512;
2512: estado = 2513;
2513: estado = 2514;
2514: estado = 2515;
2515: estado = 2516;
2516: estado = 2517;
2517: estado = 2518;
2518: estado = 2519;
2519: estado = 2520;
2520: estado = 2521;
2521: estado = 2522;
2522: estado = 2523;
2523: estado = 2524;
2524: estado = 2525;
2525: estado = 2526;
2526: estado = 2527;
2527: estado = 2528;
2528: estado = 2529;
2529: estado = 2530;
2530: estado = 2531;
2531: estado = 2532;
2532: estado = 2533;
2533: estado = 2534;
2534: estado = 2535;
2535: estado = 2536;
2536: estado = 2537;
2537: estado = 2538;
2538: estado = 2539;
2539: estado = 2540;
2540: estado = 2541;
2541: estado = 2542;
2542: estado = 2543;
2543: estado = 2544;
2544: estado = 2545;
2545: estado = 2546;
2546: estado = 2547;
2547: estado = 2548;
2548: estado = 2549;
2549: estado = 2550;
2550: estado = 2551;
2551: estado = 2552;
2552: estado = 2553;
2553: estado = 2554;
2554: estado = 2555;
2555: estado = 2556;
2556: estado = 2557;
2557: estado = 2558;
2558: estado = 2559;
2559: estado = 2560;
2560: estado = 2561;
2561: estado = 2562;
2562: estado = 2563;
2563: estado = 2564;
2564: estado = 2565;
2565: estado = 2566;
2566: estado = 2567;
2567: estado = 2568;
2568: estado = 2569;
2569: estado = 2570;
2570: estado = 2571;
2571: estado = 2572;
2572: estado = 2573;
2573: estado = 2574;
2574: estado = 2575;
2575: estado = 2576;
2576: estado = 2577;
2577: estado = 2578;
2578: estado = 2579;
2579: estado = 2580;
2580: estado = 2581;
2581: estado = 2582;
2582: estado = 2583;
2583: estado = 2584;
2584: estado = 2585;
2585: estado = 2586;
2586: estado = 2587;
2587: estado = 2588;
2588: estado = 2589;
2589: estado = 2590;
2590: estado = 2591;
2591: estado = 2592;
2592: estado = 2593;
2593: estado = 2594;
2594: estado = 2595;
2595: estado = 2596;
2596: estado = 2597;
2597: estado = 2598;
2598: estado = 2599;
2599: estado = 2600;
2600: estado = 2601;
2601: estado = 2602;
2602: estado = 2603;
2603: estado = 2604;
2604: estado = 2605;
2605: estado = 2606;
2606: estado = 2607;
2607: estado = 2608;
2608: estado = 2609;
2609: estado = 2610;
2610: estado = 2611;
2611: estado = 2612;
2612: estado = 2613;
2613: estado = 2614;
2614: estado = 2615;
2615: estado = 2616;
2616: estado = 2617;
2617: estado = 2618;
2618: estado = 2619;
2619: estado = 2620;
2620: estado = 2621;
2621: estado = 2622;
2622: estado = 2623;
2623: estado = 2624;
2624: estado = 2625;
2625: estado = 2626;
2626: estado = 2627;
2627: estado = 2628;
2628: estado = 2629;
2629: estado = 2630;
2630: estado = 2631;
2631: estado = 2632;
2632: estado = 2633;
2633: estado = 2634;
2634: estado = 2635;
2635: estado = 2636;
2636: estado = 2637;
2637: estado = 2638;
2638: estado = 2639;
2639: estado = 2640;
2640: estado = 2641;
2641: estado = 2642;
2642: estado = 2643;
2643: estado = 2644;
2644: estado = 2645;
2645: estado = 2646;
2646: estado = 2647;
2647: estado = 2648;
2648: estado = 2649;
2649: estado = 2650;
2650: estado = 2651;
2651: estado = 2652;
2652: estado = 2653;
2653: estado = 2654;
2654: estado = 2655;
2655: estado = 2656;
2656: estado = 2657;
2657: estado = 2658;
2658: estado = 2659;
2659: estado = 2660;
2660: estado = 2661;
2661: estado = 2662;
2662: estado = 2663;
2663: estado = 2664;
2664: estado = 2665;
2665: estado = 2666;
2666: estado = 2667;
2667: estado = 2668;
2668: estado = 2669;
2669: estado = 2670;
2670: estado = 2671;
2671: estado = 2672;
2672: estado = 2673;
2673: estado = 2674;
2674: estado = 2675;
2675: estado = 2676;
2676: estado = 2677;
2677: estado = 2678;
2678: estado = 2679;
2679: estado = 2680;
2680: estado = 2681;
2681: estado = 2682;
2682: estado = 2683;
2683: estado = 2684;
2684: estado = 2685;
2685: estado = 2686;
2686: estado = 2687;
2687: estado = 2688;
2688: estado = 2689;
2689: estado = 2690;
2690: estado = 2691;
2691: estado = 2692;
2692: estado = 2693;
2693: estado = 2694;
2694: estado = 2695;
2695: estado = 2696;
2696: estado = 2697;
2697: estado = 2698;
2698: estado = 2699;
2699: estado = 2700;
2700: estado = 2701;
2701: estado = 2702;
2702: estado = 2703;
2703: estado = 2704;
2704: estado = 2705;
2705: estado = 2706;
2706: estado = 2707;
2707: estado = 2708;
2708: estado = 2709;
2709: estado = 2710;
2710: estado = 2711;
2711: estado = 2712;
2712: estado = 2713;
2713: estado = 2714;
2714: estado = 2715;
2715: estado = 2716;
2716: estado = 2717;
2717: estado = 2718;
2718: estado = 2719;
2719: estado = 2720;
2720: estado = 2721;
2721: estado = 2722;
2722: estado = 2723;
2723: estado = 2724;
2724: estado = 2725;
2725: estado = 2726;
2726: estado = 2727;
2727: estado = 2728;
2728: estado = 2729;
2729: estado = 2730;
2730: estado = 2731;
2731: estado = 2732;
2732: estado = 2733;
2733: estado = 2734;
2734: estado = 2735;
2735: estado = 2736;
2736: estado = 2737;
2737: estado = 2738;
2738: estado = 2739;
2739: estado = 2740;
2740: estado = 2741;
2741: estado = 2742;
2742: estado = 2743;
2743: estado = 2744;
2744: estado = 2745;
2745: estado = 2746;
2746: estado = 2747;
2747: estado = 2748;
2748: estado = 2749;
2749: estado = 2750;
2750: estado = 2751;
2751: estado = 2752;
2752: estado = 2753;
2753: estado = 2754;
2754: estado = 2755;
2755: estado = 2756;
2756: estado = 2757;
2757: estado = 2758;
2758: estado = 2759;
2759: estado = 2760;
2760: estado = 2761;
2761: estado = 2762;
2762: estado = 2763;
2763: estado = 2764;
2764: estado = 2765;
2765: estado = 2766;
2766: estado = 2767;
2767: estado = 2768;
2768: estado = 2769;
2769: estado = 2770;
2770: estado = 2771;
2771: estado = 2772;
2772: estado = 2773;
2773: estado = 2774;
2774: estado = 2775;
2775: estado = 2776;
2776: estado = 2777;
2777: estado = 2778;
2778: estado = 2779;
2779: estado = 2780;
2780: estado = 2781;
2781: estado = 2782;
2782: estado = 2783;
2783: estado = 2784;
2784: estado = 2785;
2785: estado = 2786;
2786: estado = 2787;
2787: estado = 2788;
2788: estado = 2789;
2789: estado = 2790;
2790: estado = 2791;
2791: estado = 2792;
2792: estado = 2793;
2793: estado = 2794;
2794: estado = 2795;
2795: estado = 2796;
2796: estado = 2797;
2797: estado = 2798;
2798: estado = 2799;
2799: estado = 2800;
2800: estado = 2801;
2801: estado = 2802;
2802: estado = 2803;
2803: estado = 2804;
2804: estado = 2805;
2805: estado = 2806;
2806: estado = 2807;
2807: estado = 2808;
2808: estado = 2809;
2809: estado = 2810;
2810: estado = 2811;
2811: estado = 2812;
2812: estado = 2813;
2813: estado = 2814;
2814: estado = 2815;
2815: estado = 2816;
2816: estado = 2817;
2817: estado = 2818;
2818: estado = 2819;
2819: estado = 2820;
2820: estado = 2821;
2821: estado = 2822;
2822: estado = 2823;
2823: estado = 2824;
2824: estado = 2825;
2825: estado = 2826;
2826: estado = 2827;
2827: estado = 2828;
2828: estado = 2829;
2829: estado = 2830;
2830: estado = 2831;
2831: estado = 2832;
2832: estado = 2833;
2833: estado = 2834;
2834: estado = 2835;
2835: estado = 2836;
2836: estado = 2837;
2837: estado = 2838;
2838: estado = 2839;
2839: estado = 2840;
2840: estado = 2841;
2841: estado = 2842;
2842: estado = 2843;
2843: estado = 2844;
2844: estado = 2845;
2845: estado = 2846;
2846: estado = 2847;
2847: estado = 2848;
2848: estado = 2849;
2849: estado = 2850;
2850: estado = 2851;
2851: estado = 2852;
2852: estado = 2853;
2853: estado = 2854;
2854: estado = 2855;
2855: estado = 2856;
2856: estado = 2857;
2857: estado = 2858;
2858: estado = 2859;
2859: estado = 2860;
2860: estado = 2861;
2861: estado = 2862;
2862: estado = 2863;
2863: estado = 2864;
2864: estado = 2865;
2865: estado = 2866;
2866: estado = 2867;
2867: estado = 2868;
2868: estado = 2869;
2869: estado = 2870;
2870: estado = 2871;
2871: estado = 2872;
2872: estado = 2873;
2873: estado = 2874;
2874: estado = 2875;
2875: estado = 2876;
2876: estado = 2877;
2877: estado = 2878;
2878: estado = 2879;
2879: estado = 2880;
2880: estado = 2881;
2881: estado = 2882;
2882: estado = 2883;
2883: estado = 2884;
2884: estado = 2885;
2885: estado = 2886;
2886: estado = 2887;
2887: estado = 2888;
2888: estado = 2889;
2889: estado = 2890;
2890: estado = 2891;
2891: estado = 2892;
2892: estado = 2893;
2893: estado = 2894;
2894: estado = 2895;
2895: estado = 2896;
2896: estado = 2897;
2897: estado = 2898;
2898: estado = 2899;
2899: estado = 2900;
2900: estado = 2901;
2901: estado = 2902;
2902: estado = 2903;
2903: estado = 2904;
2904: estado = 2905;
2905: estado = 2906;
2906: estado = 2907;
2907: estado = 2908;
2908: estado = 2909;
2909: estado = 2910;
2910: estado = 2911;
2911: estado = 2912;
2912: estado = 2913;
2913: estado = 2914;
2914: estado = 2915;
2915: estado = 2916;
2916: estado = 2917;
2917: estado = 2918;
2918: estado = 2919;
2919: estado = 2920;
2920: estado = 2921;
2921: estado = 2922;
2922: estado = 2923;
2923: estado = 2924;
2924: estado = 2925;
2925: estado = 2926;
2926: estado = 2927;
2927: estado = 2928;
2928: estado = 2929;
2929: estado = 2930;
2930: estado = 2931;
2931: estado = 2932;
2932: estado = 2933;
2933: estado = 2934;
2934: estado = 2935;
2935: estado = 2936;
2936: estado = 2937;
2937: estado = 2938;
2938: estado = 2939;
2939: estado = 2940;
2940: estado = 2941;
2941: estado = 2942;
2942: estado = 2943;
2943: estado = 2944;
2944: estado = 2945;
2945: estado = 2946;
2946: estado = 2947;
2947: estado = 2948;
2948: estado = 2949;
2949: estado = 2950;
2950: estado = 2951;
2951: estado = 2952;
2952: estado = 2953;
2953: estado = 2954;
2954: estado = 2955;
2955: estado = 2956;
2956: estado = 2957;
2957: estado = 2958;
2958: estado = 2959;
2959: estado = 2960;
2960: estado = 2961;
2961: estado = 2962;
2962: estado = 2963;
2963: estado = 2964;
2964: estado = 2965;
2965: estado = 2966;
2966: estado = 2967;
2967: estado = 2968;
2968: estado = 2969;
2969: estado = 2970;
2970: estado = 2971;
2971: estado = 2972;
2972: estado = 2973;
2973: estado = 2974;
2974: estado = 2975;
2975: estado = 2976;
2976: estado = 2977;
2977: estado = 2978;
2978: estado = 2979;
2979: estado = 2980;
2980: estado = 2981;
2981: estado = 2982;
2982: estado = 2983;
2983: estado = 2984;
2984: estado = 2985;
2985: estado = 2986;
2986: estado = 2987;
2987: estado = 2988;
2988: estado = 2989;
2989: estado = 2990;
2990: estado = 2991;
2991: estado = 2992;
2992: estado = 2993;
2993: estado = 2994;
2994: estado = 2995;
2995: estado = 2996;
2996: estado = 2997;
2997: estado = 2998;
2998: estado = 2999;
2999: estado = 3000;
3000: estado = 3001;
3001: estado = 3002;
3002: estado = 3003;
3003: estado = 3004;
3004: estado = 3005;
3005: estado = 3006;
3006: estado = 3007;
3007: estado = 3008;
3008: estado = 3009;
3009: estado = 3010;
3010: estado = 3011;
3011: estado = 3012;
3012: estado = 3013;
3013: estado = 3014;
3014: estado = 3015;
3015: estado = 3016;
3016: estado = 3017;
3017: estado = 3018;
3018: estado = 3019;
3019: estado = 3020;
3020: estado = 3021;
3021: estado = 3022;
3022: estado = 3023;
3023: estado = 3024;
3024: estado = 3025;
3025: estado = 3026;
3026: estado = 3027;
3027: estado = 3028;
3028: estado = 3029;
3029: estado = 3030;
3030: estado = 3031;
3031: estado = 3032;
3032: estado = 3033;
3033: estado = 3034;
3034: estado = 3035;
3035: estado = 3036;
3036: estado = 3037;
3037: estado = 3038;
3038: estado = 3039;
3039: estado = 3040;
3040: estado = 3041;
3041: estado = 3042;
3042: estado = 3043;
3043: estado = 3044;
3044: estado = 3045;
3045: estado = 3046;
3046: estado = 3047;
3047: estado = 3048;
3048: estado = 3049;
3049: estado = 3050;
3050: estado = 3051;
3051: estado = 3052;
3052: estado = 3053;
3053: estado = 3054;
3054: estado = 3055;
3055: estado = 3056;
3056: estado = 3057;
3057: estado = 3058;
3058: estado = 3059;
3059: estado = 3060;
3060: estado = 3061;
3061: estado = 3062;
3062: estado = 3063;
3063: estado = 3064;
3064: estado = 3065;
3065: estado = 3066;
3066: estado = 3067;
3067: estado = 3068;
3068: estado = 3069;
3069: estado = 3070;
3070: estado = 3071;
3071: estado = 3072;
3072: estado = 3073;
3073: estado = 3074;
3074: estado = 3075;
3075: estado = 3076;
3076: estado = 3077;
3077: estado = 3078;
3078: estado = 3079;
3079: estado = 3080;
3080: estado = 3081;
3081: estado = 3082;
3082: estado = 3083;
3083: estado = 3084;
3084: estado = 3085;
3085: estado = 3086;
3086: estado = 3087;
3087: estado = 3088;
3088: estado = 3089;
3089: estado = 3090;
3090: estado = 3091;
3091: estado = 3092;
3092: estado = 3093;
3093: estado = 3094;
3094: estado = 3095;
3095: estado = 3096;
3096: estado = 3097;
3097: estado = 3098;
3098: estado = 3099;
3099: estado = 3100;
3100: estado = 3101;
3101: estado = 3102;
3102: estado = 3103;
3103: estado = 3104;
3104: estado = 3105;
3105: estado = 3106;
3106: estado = 3107;
3107: estado = 3108;
3108: estado = 3109;
3109: estado = 3110;
3110: estado = 3111;
3111: estado = 3112;
3112: estado = 3113;
3113: estado = 3114;
3114: estado = 3115;
3115: estado = 3116;
3116: estado = 3117;
3117: estado = 3118;
3118: estado = 3119;
3119: estado = 3120;
3120: estado = 3121;
3121: estado = 3122;
3122: estado = 3123;
3123: estado = 3124;
3124: estado = 3125;
3125: estado = 3126;
3126: estado = 3127;
3127: estado = 3128;
3128: estado = 3129;
3129: estado = 3130;
3130: estado = 3131;
3131: estado = 3132;
3132: estado = 3133;
3133: estado = 3134;
3134: estado = 3135;
3135: estado = 3136;
3136: estado = 3137;
3137: estado = 3138;
3138: estado = 3139;
3139: estado = 3140;
3140: estado = 3141;
3141: estado = 3142;
3142: estado = 3143;
3143: estado = 3144;
3144: estado = 3145;
3145: estado = 3146;
3146: estado = 3147;
3147: estado = 3148;
3148: estado = 3149;
3149: estado = 3150;
3150: estado = 3151;
3151: estado = 3152;
3152: estado = 3153;
3153: estado = 3154;
3154: estado = 3155;
3155: estado = 3156;
3156: estado = 3157;
3157: estado = 3158;
3158: estado = 3159;
3159: estado = 3160;
3160: estado = 3161;
3161: estado = 3162;
3162: estado = 3163;
3163: estado = 3164;
3164: estado = 3165;
3165: estado = 3166;
3166: estado = 3167;
3167: estado = 3168;
3168: estado = 3169;
3169: estado = 3170;
3170: estado = 3171;
3171: estado = 3172;
3172: estado = 3173;
3173: estado = 3174;
3174: estado = 3175;
3175: estado = 3176;
3176: estado = 3177;
3177: estado = 3178;
3178: estado = 3179;
3179: estado = 3180;
3180: estado = 3181;
3181: estado = 3182;
3182: estado = 3183;
3183: estado = 3184;
3184: estado = 3185;
3185: estado = 3186;
3186: estado = 3187;
3187: estado = 3188;
3188: estado = 3189;
3189: estado = 3190;
3190: estado = 3191;
3191: estado = 3192;
3192: estado = 3193;
3193: estado = 3194;
3194: estado = 3195;
3195: estado = 3196;
3196: estado = 3197;
3197: estado = 3198;
3198: estado = 3199;
3199: estado = 3200;
3200: estado = 3201;
3201: estado = 3202;
3202: estado = 3203;
3203: estado = 3204;
3204: estado = 3205;
3205: estado = 3206;
3206: estado = 3207;
3207: estado = 3208;
3208: estado = 3209;
3209: estado = 3210;
3210: estado = 3211;
3211: estado = 3212;
3212: estado = 3213;
3213: estado = 3214;
3214: estado = 3215;
3215: estado = 3216;
3216: estado = 3217;
3217: estado = 3218;
3218: estado = 3219;
3219: estado = 3220;
3220: estado = 3221;
3221: estado = 3222;
3222: estado = 3223;
3223: estado = 3224;
3224: estado = 3225;
3225: estado = 3226;
3226: estado = 3227;
3227: estado = 3228;
3228: estado = 3229;
3229: estado = 3230;
3230: estado = 3231;
3231: estado = 3232;
3232: estado = 3233;
3233: estado = 3234;
3234: estado = 3235;
3235: estado = 3236;
3236: estado = 3237;
3237: estado = 3238;
3238: estado = 3239;
3239: estado = 3240;
3240: estado = 3241;
3241: estado = 3242;
3242: estado = 3243;
3243: estado = 3244;
3244: estado = 3245;
3245: estado = 3246;
3246: estado = 3247;
3247: estado = 3248;
3248: estado = 3249;
3249: estado = 3250;
3250: estado = 3251;
3251: estado = 3252;
3252: estado = 3253;
3253: estado = 3254;
3254: estado = 3255;
3255: estado = 3256;
3256: estado = 3257;
3257: estado = 3258;
3258: estado = 3259;
3259: estado = 3260;
3260: estado = 3261;
3261: estado = 3262;
3262: estado = 3263;
3263: estado = 3264;
3264: estado = 3265;
3265: estado = 3266;
3266: estado = 3267;
3267: estado = 3268;
3268: estado = 3269;
3269: estado = 3270;
3270: estado = 3271;
3271: estado = 3272;
3272: estado = 3273;
3273: estado = 3274;
3274: estado = 3275;
3275: estado = 3276;
3276: estado = 3277;
3277: estado = 3278;
3278: estado = 3279;
3279: estado = 3280;
3280: estado = 3281;
3281: estado = 3282;
3282: estado = 3283;
3283: estado = 3284;
3284: estado = 3285;
3285: estado = 3286;
3286: estado = 3287;
3287: estado = 3288;
3288: estado = 3289;
3289: estado = 3290;
3290: estado = 3291;
3291: estado = 3292;
3292: estado = 3293;
3293: estado = 3294;
3294: estado = 3295;
3295: estado = 3296;
3296: estado = 3297;
3297: estado = 3298;
3298: estado = 3299;
3299: estado = 3300;
3300: estado = 3301;
3301: estado = 3302;
3302: estado = 3303;
3303: estado = 3304;
3304: estado = 3305;
3305: estado = 3306;
3306: estado = 3307;
3307: estado = 3308;
3308: estado = 3309;
3309: estado = 3310;
3310: estado = 3311;
3311: estado = 3312;
3312: estado = 3313;
3313: estado = 3314;
3314: estado = 3315;
3315: estado = 3316;
3316: estado = 3317;
3317: estado = 3318;
3318: estado = 3319;
3319: estado = 3320;
3320: estado = 3321;
3321: estado = 3322;
3322: estado = 3323;
3323: estado = 3324;
3324: estado = 3325;
3325: estado = 3326;
3326: estado = 3327;
3327: estado = 3328;
3328: estado = 3329;
3329: estado = 3330;
3330: estado = 3331;
3331: estado = 3332;
3332: estado = 3333;
3333: estado = 3334;
3334: estado = 3335;
3335: estado = 3336;
3336: estado = 3337;
3337: estado = 3338;
3338: estado = 3339;
3339: estado = 3340;
3340: estado = 3341;
3341: estado = 3342;
3342: estado = 3343;
3343: estado = 3344;
3344: estado = 3345;
3345: estado = 3346;
3346: estado = 3347;
3347: estado = 3348;
3348: estado = 3349;
3349: estado = 3350;
3350: estado = 3351;
3351: estado = 3352;
3352: estado = 3353;
3353: estado = 3354;
3354: estado = 3355;
3355: estado = 3356;
3356: estado = 3357;
3357: estado = 3358;
3358: estado = 3359;
3359: estado = 3360;
3360: estado = 3361;
3361: estado = 3362;
3362: estado = 3363;
3363: estado = 3364;
3364: estado = 3365;
3365: estado = 3366;
3366: estado = 3367;
3367: estado = 3368;
3368: estado = 3369;
3369: estado = 3370;
3370: estado = 3371;
3371: estado = 3372;
3372: estado = 3373;
3373: estado = 3374;
3374: estado = 3375;
3375: estado = 3376;
3376: estado = 3377;
3377: estado = 3378;
3378: estado = 3379;
3379: estado = 3380;
3380: estado = 3381;
3381: estado = 3382;
3382: estado = 3383;
3383: estado = 3384;
3384: estado = 3385;
3385: estado = 3386;
3386: estado = 3387;
3387: estado = 3388;
3388: estado = 3389;
3389: estado = 3390;
3390: estado = 3391;
3391: estado = 3392;
3392: estado = 3393;
3393: estado = 3394;
3394: estado = 3395;
3395: estado = 3396;
3396: estado = 3397;
3397: estado = 3398;
3398: estado = 3399;
3399: estado = 3400;
3400: estado = 3401;
3401: estado = 3402;
3402: estado = 3403;
3403: estado = 3404;
3404: estado = 3405;
3405: estado = 3406;
3406: estado = 3407;
3407: estado = 3408;
3408: estado = 3409;
3409: estado = 3410;
3410: estado = 3411;
3411: estado = 3412;
3412: estado = 3413;
3413: estado = 3414;
3414: estado = 3415;
3415: estado = 3416;
3416: estado = 3417;
3417: estado = 3418;
3418: estado = 3419;
3419: estado = 3420;
3420: estado = 3421;
3421: estado = 3422;
3422: estado = 3423;
3423: estado = 3424;
3424: estado = 3425;
3425: estado = 3426;
3426: estado = 3427;
3427: estado = 3428;
3428: estado = 3429;
3429: estado = 3430;
3430: estado = 3431;
3431: estado = 3432;
3432: estado = 3433;
3433: estado = 3434;
3434: estado = 3435;
3435: estado = 3436;
3436: estado = 3437;
3437: estado = 3438;
3438: estado = 3439;
3439: estado = 3440;
3440: estado = 3441;
3441: estado = 3442;
3442: estado = 3443;
3443: estado = 3444;
3444: estado = 3445;
3445: estado = 3446;
3446: estado = 3447;
3447: estado = 3448;
3448: estado = 3449;
3449: estado = 3450;
3450: estado = 3451;
3451: estado = 3452;
3452: estado = 3453;
3453: estado = 3454;
3454: estado = 3455;
3455: estado = 3456;
3456: estado = 3457;
3457: estado = 3458;
3458: estado = 3459;
3459: estado = 3460;
3460: estado = 3461;
3461: estado = 3462;
3462: estado = 3463;
3463: estado = 3464;
3464: estado = 3465;
3465: estado = 3466;
3466: estado = 3467;
3467: estado = 3468;
3468: estado = 3469;
3469: estado = 3470;
3470: estado = 3471;
3471: estado = 3472;
3472: estado = 3473;
3473: estado = 3474;
3474: estado = 3475;
3475: estado = 3476;
3476: estado = 3477;
3477: estado = 3478;
3478: estado = 3479;
3479: estado = 3480;
3480: estado = 3481;
3481: estado = 3482;
3482: estado = 3483;
3483: estado = 3484;
3484: estado = 3485;
3485: estado = 3486;
3486: estado = 3487;
3487: estado = 3488;
3488: estado = 3489;
3489: estado = 3490;
3490: estado = 3491;
3491: estado = 3492;
3492: estado = 3493;
3493: estado = 3494;
3494: estado = 3495;
3495: estado = 3496;
3496: estado = 3497;
3497: estado = 3498;
3498: estado = 3499;
3499: estado = 3500;
3500: estado = 3501;
3501: estado = 3502;
3502: estado = 3503;
3503: estado = 3504;
3504: estado = 3505;
3505: estado = 3506;
3506: estado = 3507;
3507: estado = 3508;
3508: estado = 3509;
3509: estado = 3510;
3510: estado = 3511;
3511: estado = 3512;
3512: estado = 3513;
3513: estado = 3514;
3514: estado = 3515;
3515: estado = 3516;
3516: estado = 3517;
3517: estado = 3518;
3518: estado = 3519;
3519: estado = 3520;
3520: estado = 3521;
3521: estado = 3522;
3522: estado = 3523;
3523: estado = 3524;
3524: estado = 3525;
3525: estado = 3526;
3526: estado = 3527;
3527: estado = 3528;
3528: estado = 3529;
3529: estado = 3530;
3530: estado = 3531;
3531: estado = 3532;
3532: estado = 3533;
3533: estado = 3534;
3534: estado = 3535;
3535: estado = 3536;
3536: estado = 3537;
3537: estado = 3538;
3538: estado = 3539;
3539: estado = 3540;
3540: estado = 3541;
3541: estado = 3542;
3542: estado = 3543;
3543: estado = 3544;
3544: estado = 3545;
3545: estado = 3546;
3546: estado = 3547;
3547: estado = 3548;
3548: estado = 3549;
3549: estado = 3550;
3550: estado = 3551;
3551: estado = 3552;
3552: estado = 3553;
3553: estado = 3554;
3554: estado = 3555;
3555: estado = 3556;
3556: estado = 3557;
3557: estado = 3558;
3558: estado = 3559;
3559: estado = 3560;
3560: estado = 3561;
3561: estado = 3562;
3562: estado = 3563;
3563: estado = 3564;
3564: estado = 3565;
3565: estado = 3566;
3566: estado = 3567;
3567: estado = 3568;
3568: estado = 3569;
3569: estado = 3570;
3570: estado = 3571;
3571: estado = 3572;
3572: estado = 3573;
3573: estado = 3574;
3574: estado = 3575;
3575: estado = 3576;
3576: estado = 3577;
3577: estado = 3578;
3578: estado = 3579;
3579: estado = 3580;
3580: estado = 3581;
3581: estado = 3582;
3582: estado = 3583;
3583: estado = 3584;
3584: estado = 3585;
3585: estado = 3586;
3586: estado = 3587;
3587: estado = 3588;
3588: estado = 3589;
3589: estado = 3590;
3590: estado = 3591;
3591: estado = 3592;
3592: estado = 3593;
3593: estado = 3594;
3594: estado = 3595;
3595: estado = 3596;
3596: estado = 3597;
3597: estado = 3598;
3598: estado = 3599;
3599: estado = 3600;
3600: estado = 3601;
3601: estado = 3602;
3602: estado = 3603;
3603: estado = 3604;
3604: estado = 3605;
3605: estado = 3606;
3606: estado = 3607;
3607: estado = 3608;
3608: estado = 3609;
3609: estado = 3610;
3610: estado = 3611;
3611: estado = 3612;
3612: estado = 3613;
3613: estado = 3614;
3614: estado = 3615;
3615: estado = 3616;
3616: estado = 3617;
3617: estado = 3618;
3618: estado = 3619;
3619: estado = 3620;
3620: estado = 3621;
3621: estado = 3622;
3622: estado = 3623;
3623: estado = 3624;
3624: estado = 3625;
3625: estado = 3626;
3626: estado = 3627;
3627: estado = 3628;
3628: estado = 3629;
3629: estado = 3630;
3630: estado = 3631;
3631: estado = 3632;
3632: estado = 3633;
3633: estado = 3634;
3634: estado = 3635;
3635: estado = 3636;
3636: estado = 3637;
3637: estado = 3638;
3638: estado = 3639;
3639: estado = 3640;
3640: estado = 3641;
3641: estado = 3642;
3642: estado = 3643;
3643: estado = 3644;
3644: estado = 3645;
3645: estado = 3646;
3646: estado = 3647;
3647: estado = 3648;
3648: estado = 3649;
3649: estado = 3650;
3650: estado = 3651;
3651: estado = 3652;
3652: estado = 3653;
3653: estado = 3654;
3654: estado = 3655;
3655: estado = 3656;
3656: estado = 3657;
3657: estado = 3658;
3658: estado = 3659;
3659: estado = 3660;
3660: estado = 3661;
3661: estado = 3662;
3662: estado = 3663;
3663: estado = 3664;
3664: estado = 3665;
3665: estado = 3666;
3666: estado = 3667;
3667: estado = 3668;
3668: estado = 3669;
3669: estado = 3670;
3670: estado = 3671;
3671: estado = 3672;
3672: estado = 3673;
3673: estado = 3674;
3674: estado = 3675;
3675: estado = 3676;
3676: estado = 3677;
3677: estado = 3678;
3678: estado = 3679;
3679: estado = 3680;
3680: estado = 3681;
3681: estado = 3682;
3682: estado = 3683;
3683: estado = 3684;
3684: estado = 3685;
3685: estado = 3686;
3686: estado = 3687;
3687: estado = 3688;
3688: estado = 3689;
3689: estado = 3690;
3690: estado = 3691;
3691: estado = 3692;
3692: estado = 3693;
3693: estado = 3694;
3694: estado = 3695;
3695: estado = 3696;
3696: estado = 3697;
3697: estado = 3698;
3698: estado = 3699;
3699: estado = 3700;
3700: estado = 3701;
3701: estado = 3702;
3702: estado = 3703;
3703: estado = 3704;
3704: estado = 3705;
3705: estado = 3706;
3706: estado = 3707;
3707: estado = 3708;
3708: estado = 3709;
3709: estado = 3710;
3710: estado = 3711;
3711: estado = 3712;
3712: estado = 3713;
3713: estado = 3714;
3714: estado = 3715;
3715: estado = 3716;
3716: estado = 3717;
3717: estado = 3718;
3718: estado = 3719;
3719: estado = 3720;
3720: estado = 3721;
3721: estado = 3722;
3722: estado = 3723;
3723: estado = 3724;
3724: estado = 3725;
3725: estado = 3726;
3726: estado = 3727;
3727: estado = 3728;
3728: estado = 3729;
3729: estado = 3730;
3730: estado = 3731;
3731: estado = 3732;
3732: estado = 3733;
3733: estado = 3734;
3734: estado = 3735;
3735: estado = 3736;
3736: estado = 3737;
3737: estado = 3738;
3738: estado = 3739;
3739: estado = 3740;
3740: estado = 3741;
3741: estado = 3742;
3742: estado = 3743;
3743: estado = 3744;
3744: estado = 3745;
3745: estado = 3746;
3746: estado = 3747;
3747: estado = 3748;
3748: estado = 3749;
3749: estado = 3750;
3750: estado = 3751;
3751: estado = 3752;
3752: estado = 3753;
3753: estado = 3754;
3754: estado = 3755;
3755: estado = 3756;
3756: estado = 3757;
3757: estado = 3758;
3758: estado = 3759;
3759: estado = 3760;
3760: estado = 3761;
3761: estado = 3762;
3762: estado = 3763;
3763: estado = 3764;
3764: estado = 3765;
3765: estado = 3766;
3766: estado = 3767;
3767: estado = 3768;
3768: estado = 3769;
3769: estado = 3770;
3770: estado = 3771;
3771: estado = 3772;
3772: estado = 3773;
3773: estado = 3774;
3774: estado = 3775;
3775: estado = 3776;
3776: estado = 3777;
3777: estado = 3778;
3778: estado = 3779;
3779: estado = 3780;
3780: estado = 3781;
3781: estado = 3782;
3782: estado = 3783;
3783: estado = 3784;
3784: estado = 3785;
3785: estado = 3786;
3786: estado = 3787;
3787: estado = 3788;
3788: estado = 3789;
3789: estado = 3790;
3790: estado = 3791;
3791: estado = 3792;
3792: estado = 3793;
3793: estado = 3794;
3794: estado = 3795;
3795: estado = 3796;
3796: estado = 3797;
3797: estado = 3798;
3798: estado = 3799;
3799: estado = 3800;
3800: estado = 3801;
3801: estado = 3802;
3802: estado = 3803;
3803: estado = 3804;
3804: estado = 3805;
3805: estado = 3806;
3806: estado = 3807;
3807: estado = 3808;
3808: estado = 3809;
3809: estado = 3810;
3810: estado = 3811;
3811: estado = 3812;
3812: estado = 3813;
3813: estado = 3814;
3814: estado = 3815;
3815: estado = 3816;
3816: estado = 3817;
3817: estado = 3818;
3818: estado = 3819;
3819: estado = 3820;
3820: estado = 3821;
3821: estado = 3822;
3822: estado = 3823;
3823: estado = 3824;
3824: estado = 3825;
3825: estado = 3826;
3826: estado = 3827;
3827: estado = 3828;
3828: estado = 3829;
3829: estado = 3830;
3830: estado = 3831;
3831: estado = 3832;
3832: estado = 3833;
3833: estado = 3834;
3834: estado = 3835;
3835: estado = 3836;
3836: estado = 3837;
3837: estado = 3838;
3838: estado = 3839;
3839: estado = 3840;
3840: estado = 3841;
3841: estado = 3842;
3842: estado = 3843;
3843: estado = 3844;
3844: estado = 3845;
3845: estado = 3846;
3846: estado = 3847;
3847: estado = 3848;
3848: estado = 3849;
3849: estado = 3850;
3850: estado = 3851;
3851: estado = 3852;
3852: estado = 3853;
3853: estado = 3854;
3854: estado = 3855;
3855: estado = 3856;
3856: estado = 3857;
3857: estado = 3858;
3858: estado = 3859;
3859: estado = 3860;
3860: estado = 3861;
3861: estado = 3862;
3862: estado = 3863;
3863: estado = 3864;
3864: estado = 3865;
3865: estado = 3866;
3866: estado = 3867;
3867: estado = 3868;
3868: estado = 3869;
3869: estado = 3870;
3870: estado = 3871;
3871: estado = 3872;
3872: estado = 3873;
3873: estado = 3874;
3874: estado = 3875;
3875: estado = 3876;
3876: estado = 3877;
3877: estado = 3878;
3878: estado = 3879;
3879: estado = 3880;
3880: estado = 3881;
3881: estado = 3882;
3882: estado = 3883;
3883: estado = 3884;
3884: estado = 3885;
3885: estado = 3886;
3886: estado = 3887;
3887: estado = 3888;
3888: estado = 3889;
3889: estado = 3890;
3890: estado = 3891;
3891: estado = 3892;
3892: estado = 3893;
3893: estado = 3894;
3894: estado = 3895;
3895: estado = 3896;
3896: estado = 3897;
3897: estado = 3898;
3898: estado = 3899;
3899: estado = 3900;
3900: estado = 3901;
3901: estado = 3902;
3902: estado = 3903;
3903: estado = 3904;
3904: estado = 3905;
3905: estado = 3906;
3906: estado = 3907;
3907: estado = 3908;
3908: estado = 3909;
3909: estado = 3910;
3910: estado = 3911;
3911: estado = 3912;
3912: estado = 3913;
3913: estado = 3914;
3914: estado = 3915;
3915: estado = 3916;
3916: estado = 3917;
3917: estado = 3918;
3918: estado = 3919;
3919: estado = 3920;
3920: estado = 3921;
3921: estado = 3922;
3922: estado = 3923;
3923: estado = 3924;
3924: estado = 3925;
3925: estado = 3926;
3926: estado = 3927;
3927: estado = 3928;
3928: estado = 3929;
3929: estado = 3930;
3930: estado = 3931;
3931: estado = 3932;
3932: estado = 3933;
3933: estado = 3934;
3934: estado = 3935;
3935: estado = 3936;
3936: estado = 3937;
3937: estado = 3938;
3938: estado = 3939;
3939: estado = 3940;
3940: estado = 3941;
3941: estado = 3942;
3942: estado = 3943;
3943: estado = 3944;
3944: estado = 3945;
3945: estado = 3946;
3946: estado = 3947;
3947: estado = 3948;
3948: estado = 3949;
3949: estado = 3950;
3950: estado = 3951;
3951: estado = 3952;
3952: estado = 3953;
3953: estado = 3954;
3954: estado = 3955;
3955: estado = 3956;
3956: estado = 3957;
3957: estado = 3958;
3958: estado = 3959;
3959: estado = 3960;
3960: estado = 3961;
3961: estado = 3962;
3962: estado = 3963;
3963: estado = 3964;
3964: estado = 3965;
3965: estado = 3966;
3966: estado = 3967;
3967: estado = 3968;
3968: estado = 3969;
3969: estado = 3970;
3970: estado = 3971;
3971: estado = 3972;
3972: estado = 3973;
3973: estado = 3974;
3974: estado = 3975;
3975: estado = 3976;
3976: estado = 3977;
3977: estado = 3978;
3978: estado = 3979;
3979: estado = 3980;
3980: estado = 3981;
3981: estado = 3982;
3982: estado = 3983;
3983: estado = 3984;
3984: estado = 3985;
3985: estado = 3986;
3986: estado = 3987;
3987: estado = 3988;
3988: estado = 3989;
3989: estado = 3990;
3990: estado = 3991;
3991: estado = 3992;
3992: estado = 3993;
3993: estado = 3994;
3994: estado = 3995;
3995: estado = 3996;
3996: estado = 3997;
3997: estado = 3998;
3998: estado = 3999;
3999: estado = 4000;
4000: estado = 4001;
4001: estado = 4002;
4002: estado = 4003;
4003: estado = 4004;
4004: estado = 4005;
4005: estado = 4006;
4006: estado = 4007;
4007: estado = 4008;
4008: estado = 4009;
4009: estado = 4010;
4010: estado = 4011;
4011: estado = 4012;
4012: estado = 4013;
4013: estado = 4014;
4014: estado = 4015;
4015: estado = 4016;
4016: estado = 4017;
4017: estado = 4018;
4018: estado = 4019;
4019: estado = 4020;
4020: estado = 4021;
4021: estado = 4022;
4022: estado = 4023;
4023: estado = 4024;
4024: estado = 4025;
4025: estado = 4026;
4026: estado = 4027;
4027: estado = 4028;
4028: estado = 4029;
4029: estado = 4030;
4030: estado = 4031;
4031: estado = 4032;
4032: estado = 4033;
4033: estado = 4034;
4034: estado = 4035;
4035: estado = 4036;
4036: estado = 4037;
4037: estado = 4038;
4038: estado = 4039;
4039: estado = 4040;
4040: estado = 4041;
4041: estado = 4042;
4042: estado = 4043;
4043: estado = 4044;
4044: estado = 4045;
4045: estado = 4046;
4046: estado = 4047;
4047: estado = 4048;
4048: estado = 4049;
4049: estado = 4050;
4050: estado = 4051;
4051: estado = 4052;
4052: estado = 4053;
4053: estado = 4054;
4054: estado = 4055;
4055: estado = 4056;
4056: estado = 4057;
4057: estado = 4058;
4058: estado = 4059;
4059: estado = 4060;
4060: estado = 4061;
4061: estado = 4062;
4062: estado = 4063;
4063: estado = 4064;
4064: estado = 4065;
4065: estado = 4066;
4066: estado = 4067;
4067: estado = 4068;
4068: estado = 4069;
4069: estado = 4070;
4070: estado = 4071;
4071: estado = 4072;
4072: estado = 4073;
4073: estado = 4074;
4074: estado = 4075;
4075: estado = 4076;
4076: estado = 4077;
4077: estado = 4078;
4078: estado = 4079;
4079: estado = 4080;
4080: estado = 4081;
4081: estado = 4082;
4082: estado = 4083;
4083: estado = 4084;
4084: estado = 4085;
4085: estado = 4086;
4086: estado = 4087;
4087: estado = 4088;
4088: estado = 4089;
4089: estado = 4090;
4090: estado = 4091;
4091: estado = 4092;
4092: estado = 4093;
4093: estado = 4094;
4094: estado = 4095;
4095: estado = 4096;
4096: estado = 4097;
4097: estado = 4098;
4098: estado = 4099;
4099: estado = 4100;
4100: estado = 4101;
4101: estado = 4102;
4102: estado = 4103;
4103: estado = 4104;
4104: estado = 4105;
4105: estado = 4106;
4106: estado = 4107;
4107: estado = 4108;
4108: estado = 4109;
4109: estado = 4110;
4110: estado = 4111;
4111: estado = 4112;
4112: estado = 4113;
4113: estado = 4114;
4114: estado = 4115;
4115: estado = 4116;
4116: estado = 4117;
4117: estado = 4118;
4118: estado = 4119;
4119: estado = 4120;
4120: estado = 4121;
4121: estado = 4122;
4122: estado = 4123;
4123: estado = 4124;
4124: estado = 4125;
4125: estado = 4126;
4126: estado = 4127;
4127: estado = 4128;
4128: estado = 4129;
4129: estado = 4130;
4130: estado = 4131;
4131: estado = 4132;
4132: estado = 4133;
4133: estado = 4134;
4134: estado = 4135;
4135: estado = 4136;
4136: estado = 4137;
4137: estado = 4138;
4138: estado = 4139;
4139: estado = 4140;
4140: estado = 4141;
4141: estado = 4142;
4142: estado = 4143;
4143: estado = 4144;
4144: estado = 4145;
4145: estado = 4146;
4146: estado = 4147;
4147: estado = 4148;
4148: estado = 4149;
4149: estado = 4150;
4150: estado = 4151;
4151: estado = 4152;
4152: estado = 4153;
4153: estado = 4154;
4154: estado = 4155;
4155: estado = 4156;
4156: estado = 4157;
4157: estado = 4158;
4158: estado = 4159;
4159: estado = 4160;
4160: estado = 4161;
4161: estado = 4162;
4162: estado = 4163;
4163: estado = 4164;
4164: estado = 4165;
4165: estado = 4166;
4166: estado = 4167;
4167: estado = 4168;
4168: estado = 4169;
4169: estado = 4170;
4170: estado = 4171;
4171: estado = 4172;
4172: estado = 4173;
4173: estado = 4174;
4174: estado = 4175;
4175: estado = 4176;
4176: estado = 4177;
4177: estado = 4178;
4178: estado = 4179;
4179: estado = 4180;
4180: estado = 4181;
4181: estado = 4182;
4182: estado = 4183;
4183: estado = 4184;
4184: estado = 4185;
4185: estado = 4186;
4186: estado = 4187;
4187: estado = 4188;
4188: estado = 4189;
4189: estado = 4190;
4190: estado = 4191;
4191: estado = 4192;
4192: estado = 4193;
4193: estado = 4194;
4194: estado = 4195;
4195: estado = 4196;
4196: estado = 4197;
4197: estado = 4198;
4198: estado = 4199;
4199: estado = 4200;
4200: estado = 4201;
4201: estado = 4202;
4202: estado = 4203;
4203: estado = 4204;
4204: estado = 4205;
4205: estado = 4206;
4206: estado = 4207;
4207: estado = 4208;
4208: estado = 4209;
4209: estado = 4210;
4210: estado = 4211;
4211: estado = 4212;
4212: estado = 4213;
4213: estado = 4214;
4214: estado = 4215;
4215: estado = 4216;
4216: estado = 4217;
4217: estado = 4218;
4218: estado = 4219;
4219: estado = 4220;
4220: estado = 4221;
4221: estado = 4222;
4222: estado = 4223;
4223: estado = 4224;
4224: estado = 4225;
4225: estado = 4226;
4226: estado = 4227;
4227: estado = 4228;
4228: estado = 4229;
4229: estado = 4230;
4230: estado = 4231;
4231: estado = 4232;
4232: estado = 4233;
4233: estado = 4234;
4234: estado = 4235;
4235: estado = 4236;
4236: estado = 4237;
4237: estado = 4238;
4238: estado = 4239;
4239: estado = 4240;
4240: estado = 4241;
4241: estado = 4242;
4242: estado = 4243;
4243: estado = 4244;
4244: estado = 4245;
4245: estado = 4246;
4246: estado = 4247;
4247: estado = 4248;
4248: estado = 4249;
4249: estado = 4250;
4250: estado = 4251;
4251: estado = 4252;
4252: estado = 4253;
4253: estado = 4254;
4254: estado = 4255;
4255: estado = 4256;
4256: estado = 4257;
4257: estado = 4258;
4258: estado = 4259;
4259: estado = 4260;
4260: estado = 4261;
4261: estado = 4262;
4262: estado = 4263;
4263: estado = 4264;
4264: estado = 4265;
4265: estado = 4266;
4266: estado = 4267;
4267: estado = 4268;
4268: estado = 4269;
4269: estado = 4270;
4270: estado = 4271;
4271: estado = 4272;
4272: estado = 4273;
4273: estado = 4274;
4274: estado = 4275;
4275: estado = 4276;
4276: estado = 4277;
4277: estado = 4278;
4278: estado = 4279;
4279: estado = 4280;
4280: estado = 4281;
4281: estado = 4282;
4282: estado = 4283;
4283: estado = 4284;
4284: estado = 4285;
4285: estado = 4286;
4286: estado = 4287;
4287: estado = 4288;
4288: estado = 4289;
4289: estado = 4290;
4290: estado = 4291;
4291: estado = 4292;
4292: estado = 4293;
4293: estado = 4294;
4294: estado = 4295;
4295: estado = 4296;
4296: estado = 4297;
4297: estado = 4298;
4298: estado = 4299;
4299: estado = 4300;
4300: estado = 4301;
4301: estado = 4302;
4302: estado = 4303;
4303: estado = 4304;
4304: estado = 4305;
4305: estado = 4306;
4306: estado = 4307;
4307: estado = 4308;
4308: estado = 4309;
4309: estado = 4310;
4310: estado = 4311;
4311: estado = 4312;
4312: estado = 4313;
4313: estado = 4314;
4314: estado = 4315;
4315: estado = 4316;
4316: estado = 4317;
4317: estado = 4318;
4318: estado = 4319;
4319: estado = 4320;
4320: estado = 4321;
4321: estado = 4322;
4322: estado = 4323;
4323: estado = 4324;
4324: estado = 4325;
4325: estado = 4326;
4326: estado = 4327;
4327: estado = 4328;
4328: estado = 4329;
4329: estado = 4330;
4330: estado = 4331;
4331: estado = 4332;
4332: estado = 4333;
4333: estado = 4334;
4334: estado = 4335;
4335: estado = 4336;
4336: estado = 4337;
4337: estado = 4338;
4338: estado = 4339;
4339: estado = 4340;
4340: estado = 4341;
4341: estado = 4342;
4342: estado = 4343;
4343: estado = 4344;
4344: estado = 4345;
4345: estado = 4346;
4346: estado = 4347;
4347: estado = 4348;
4348: estado = 4349;
4349: estado = 4350;
4350: estado = 4351;
4351: estado = 4352;
4352: estado = 4353;
4353: estado = 4354;
4354: estado = 4355;
4355: estado = 4356;
4356: estado = 4357;
4357: estado = 4358;
4358: estado = 4359;
4359: estado = 4360;
4360: estado = 4361;
4361: estado = 4362;
4362: estado = 4363;
4363: estado = 4364;
4364: estado = 4365;
4365: estado = 4366;
4366: estado = 4367;
4367: estado = 4368;
4368: estado = 4369;
4369: estado = 4370;
4370: estado = 4371;
4371: estado = 4372;
4372: estado = 4373;
4373: estado = 4374;
4374: estado = 4375;
4375: estado = 4376;
4376: estado = 4377;
4377: estado = 4378;
4378: estado = 4379;
4379: estado = 4380;
4380: estado = 4381;
4381: estado = 4382;
4382: estado = 4383;
4383: estado = 4384;
4384: estado = 4385;
4385: estado = 4386;
4386: estado = 4387;
4387: estado = 4388;
4388: estado = 4389;
4389: estado = 4390;
4390: estado = 4391;
4391: estado = 4392;
4392: estado = 4393;
4393: estado = 4394;
4394: estado = 4395;
4395: estado = 4396;
4396: estado = 4397;
4397: estado = 4398;
4398: estado = 4399;
4399: estado = 4400;
4400: estado = 4401;
4401: estado = 4402;
4402: estado = 4403;
4403: estado = 4404;
4404: estado = 4405;
4405: estado = 4406;
4406: estado = 4407;
4407: estado = 4408;
4408: estado = 4409;
4409: estado = 4410;
4410: estado = 4411;
4411: estado = 4412;
4412: estado = 4413;
4413: estado = 4414;
4414: estado = 4415;
4415: estado = 4416;
4416: estado = 4417;
4417: estado = 4418;
4418: estado = 4419;
4419: estado = 4420;
4420: estado = 4421;
4421: estado = 4422;
4422: estado = 4423;
4423: estado = 4424;
4424: estado = 4425;
4425: estado = 4426;
4426: estado = 4427;
4427: estado = 4428;
4428: estado = 4429;
4429: estado = 4430;
4430: estado = 4431;
4431: estado = 4432;
4432: estado = 4433;
4433: estado = 4434;
4434: estado = 4435;
4435: estado = 4436;
4436: estado = 4437;
4437: estado = 4438;
4438: estado = 4439;
4439: estado = 4440;
4440: estado = 4441;
4441: estado = 4442;
4442: estado = 4443;
4443: estado = 4444;
4444: estado = 4445;
4445: estado = 4446;
4446: estado = 4447;
4447: estado = 4448;
4448: estado = 4449;
4449: estado = 4450;
4450: estado = 4451;
4451: estado = 4452;
4452: estado = 4453;
4453: estado = 4454;
4454: estado = 4455;
4455: estado = 4456;
4456: estado = 4457;
4457: estado = 4458;
4458: estado = 4459;
4459: estado = 4460;
4460: estado = 4461;
4461: estado = 4462;
4462: estado = 4463;
4463: estado = 4464;
4464: estado = 4465;
4465: estado = 4466;
4466: estado = 4467;
4467: estado = 4468;
4468: estado = 4469;
4469: estado = 4470;
4470: estado = 4471;
4471: estado = 4472;
4472: estado = 4473;
4473: estado = 4474;
4474: estado = 4475;
4475: estado = 4476;
4476: estado = 4477;
4477: estado = 4478;
4478: estado = 4479;
4479: estado = 4480;
4480: estado = 4481;
4481: estado = 4482;
4482: estado = 4483;
4483: estado = 4484;
4484: estado = 4485;
4485: estado = 4486;
4486: estado = 4487;
4487: estado = 4488;
4488: estado = 4489;
4489: estado = 4490;
4490: estado = 4491;
4491: estado = 4492;
4492: estado = 4493;
4493: estado = 4494;
4494: estado = 4495;
4495: estado = 4496;
4496: estado = 4497;
4497: estado = 4498;
4498: estado = 4499;
4499: estado = 4500;
4500: estado = 4501;
4501: estado = 4502;
4502: estado = 4503;
4503: estado = 4504;
4504: estado = 4505;
4505: estado = 4506;
4506: estado = 4507;
4507: estado = 4508;
4508: estado = 4509;
4509: estado = 4510;
4510: estado = 4511;
4511: estado = 4512;
4512: estado = 4513;
4513: estado = 4514;
4514: estado = 4515;
4515: estado = 4516;
4516: estado = 4517;
4517: estado = 4518;
4518: estado = 4519;
4519: estado = 4520;
4520: estado = 4521;
4521: estado = 4522;
4522: estado = 4523;
4523: estado = 4524;
4524: estado = 4525;
4525: estado = 4526;
4526: estado = 4527;
4527: estado = 4528;
4528: estado = 4529;
4529: estado = 4530;
4530: estado = 4531;
4531: estado = 4532;
4532: estado = 4533;
4533: estado = 4534;
4534: estado = 4535;
4535: estado = 4536;
4536: estado = 4537;
4537: estado = 4538;
4538: estado = 4539;
4539: estado = 4540;
4540: estado = 4541;
4541: estado = 4542;
4542: estado = 4543;
4543: estado = 4544;
4544: estado = 4545;
4545: estado = 4546;
4546: estado = 4547;
4547: estado = 4548;
4548: estado = 4549;
4549: estado = 4550;
4550: estado = 4551;
4551: estado = 4552;
4552: estado = 4553;
4553: estado = 4554;
4554: estado = 4555;
4555: estado = 4556;
4556: estado = 4557;
4557: estado = 4558;
4558: estado = 4559;
4559: estado = 4560;
4560: estado = 4561;
4561: estado = 4562;
4562: estado = 4563;
4563: estado = 4564;
4564: estado = 4565;
4565: estado = 4566;
4566: estado = 4567;
4567: estado = 4568;
4568: estado = 4569;
4569: estado = 4570;
4570: estado = 4571;
4571: estado = 4572;
4572: estado = 4573;
4573: estado = 4574;
4574: estado = 4575;
4575: estado = 4576;
4576: estado = 4577;
4577: estado = 4578;
4578: estado = 4579;
4579: estado = 4580;
4580: estado = 4581;
4581: estado = 4582;
4582: estado = 4583;
4583: estado = 4584;
4584: estado = 4585;
4585: estado = 4586;
4586: estado = 4587;
4587: estado = 4588;
4588: estado = 4589;
4589: estado = 4590;
4590: estado = 4591;
4591: estado = 4592;
4592: estado = 4593;
4593: estado = 4594;
4594: estado = 4595;
4595: estado = 4596;
4596: estado = 4597;
4597: estado = 4598;
4598: estado = 4599;
4599: estado = 4600;
4600: estado = 4601;
4601: estado = 4602;
4602: estado = 4603;
4603: estado = 4604;
4604: estado = 4605;
4605: estado = 4606;
4606: estado = 4607;
4607: estado = 4608;
4608: estado = 4609;
4609: estado = 4610;
4610: estado = 4611;
4611: estado = 4612;
4612: estado = 4613;
4613: estado = 4614;
4614: estado = 4615;
4615: estado = 4616;
4616: estado = 4617;
4617: estado = 4618;
4618: estado = 4619;
4619: estado = 4620;
4620: estado = 4621;
4621: estado = 4622;
4622: estado = 4623;
4623: estado = 4624;
4624: estado = 4625;
4625: estado = 4626;
4626: estado = 4627;
4627: estado = 4628;
4628: estado = 4629;
4629: estado = 4630;
4630: estado = 4631;
4631: estado = 4632;
4632: estado = 4633;
4633: estado = 4634;
4634: estado = 4635;
4635: estado = 4636;
4636: estado = 4637;
4637: estado = 4638;
4638: estado = 4639;
4639: estado = 4640;
4640: estado = 4641;
4641: estado = 4642;
4642: estado = 4643;
4643: estado = 4644;
4644: estado = 4645;
4645: estado = 4646;
4646: estado = 4647;
4647: estado = 4648;
4648: estado = 4649;
4649: estado = 4650;
4650: estado = 4651;
4651: estado = 4652;
4652: estado = 4653;
4653: estado = 4654;
4654: estado = 4655;
4655: estado = 4656;
4656: estado = 4657;
4657: estado = 4658;
4658: estado = 4659;
4659: estado = 4660;
4660: estado = 4661;
4661: estado = 4662;
4662: estado = 4663;
4663: estado = 4664;
4664: estado = 4665;
4665: estado = 4666;
4666: estado = 4667;
4667: estado = 4668;
4668: estado = 4669;
4669: estado = 4670;
4670: estado = 4671;
4671: estado = 4672;
4672: estado = 4673;
4673: estado = 4674;
4674: estado = 4675;
4675: estado = 4676;
4676: estado = 4677;
4677: estado = 4678;
4678: estado = 4679;
4679: estado = 4680;
4680: estado = 4681;
4681: estado = 4682;
4682: estado = 4683;
4683: estado = 4684;
4684: estado = 4685;
4685: estado = 4686;
4686: estado = 4687;
4687: estado = 4688;
4688: estado = 4689;
4689: estado = 4690;
4690: estado = 4691;
4691: estado = 4692;
4692: estado = 4693;
4693: estado = 4694;
4694: estado = 4695;
4695: estado = 4696;
4696: estado = 4697;
4697: estado = 4698;
4698: estado = 4699;
4699: estado = 4700;
4700: estado = 4701;
4701: estado = 4702;
4702: estado = 4703;
4703: estado = 4704;
4704: estado = 4705;
4705: estado = 4706;
4706: estado = 4707;
4707: estado = 4708;
4708: estado = 4709;
4709: estado = 4710;
4710: estado = 4711;
4711: estado = 4712;
4712: estado = 4713;
4713: estado = 4714;
4714: estado = 4715;
4715: estado = 4716;
4716: estado = 4717;
4717: estado = 4718;
4718: estado = 4719;
4719: estado = 4720;
4720: estado = 4721;
4721: estado = 4722;
4722: estado = 4723;
4723: estado = 4724;
4724: estado = 4725;
4725: estado = 4726;
4726: estado = 4727;
4727: estado = 4728;
4728: estado = 4729;
4729: estado = 4730;
4730: estado = 4731;
4731: estado = 4732;
4732: estado = 4733;
4733: estado = 4734;
4734: estado = 4735;
4735: estado = 4736;
4736: estado = 4737;
4737: estado = 4738;
4738: estado = 4739;
4739: estado = 4740;
4740: estado = 4741;
4741: estado = 4742;
4742: estado = 4743;
4743: estado = 4744;
4744: estado = 4745;
4745: estado = 4746;
4746: estado = 4747;
4747: estado = 4748;
4748: estado = 4749;
4749: estado = 4750;
4750: estado = 4751;
4751: estado = 4752;
4752: estado = 4753;
4753: estado = 4754;
4754: estado = 4755;
4755: estado = 4756;
4756: estado = 4757;
4757: estado = 4758;
4758: estado = 4759;
4759: estado = 4760;
4760: estado = 4761;
4761: estado = 4762;
4762: estado = 4763;
4763: estado = 4764;
4764: estado = 4765;
4765: estado = 4766;
4766: estado = 4767;
4767: estado = 4768;
4768: estado = 4769;
4769: estado = 4770;
4770: estado = 4771;
4771: estado = 4772;
4772: estado = 4773;
4773: estado = 4774;
4774: estado = 4775;
4775: estado = 4776;
4776: estado = 4777;
4777: estado = 4778;
4778: estado = 4779;
4779: estado = 4780;
4780: estado = 4781;
4781: estado = 4782;
4782: estado = 4783;
4783: estado = 4784;
4784: estado = 4785;
4785: estado = 4786;
4786: estado = 4787;
4787: estado = 4788;
4788: estado = 4789;
4789: estado = 4790;
4790: estado = 4791;
4791: estado = 4792;
4792: estado = 4793;
4793: estado = 4794;
4794: estado = 4795;
4795: estado = 4796;
4796: estado = 4797;
4797: estado = 4798;
4798: estado = 4799;
4799: estado = 4800;
4800: estado = 4801;
4801: estado = 4802;
4802: estado = 4803;
4803: estado = 4804;
4804: estado = 4805;
4805: estado = 4806;
4806: estado = 4807;
4807: estado = 4808;
4808: estado = 4809;
4809: estado = 4810;
4810: estado = 4811;
4811: estado = 4812;
4812: estado = 4813;
4813: estado = 4814;
4814: estado = 4815;
4815: estado = 4816;
4816: estado = 4817;
4817: estado = 4818;
4818: estado = 4819;
4819: estado = 4820;
4820: estado = 4821;
4821: estado = 4822;
4822: estado = 4823;
4823: estado = 4824;
4824: estado = 4825;
4825: estado = 4826;
4826: estado = 4827;
4827: estado = 4828;
4828: estado = 4829;
4829: estado = 4830;
4830: estado = 4831;
4831: estado = 4832;
4832: estado = 4833;
4833: estado = 4834;
4834: estado = 4835;
4835: estado = 4836;
4836: estado = 4837;
4837: estado = 4838;
4838: estado = 4839;
4839: estado = 4840;
4840: estado = 4841;
4841: estado = 4842;
4842: estado = 4843;
4843: estado = 4844;
4844: estado = 4845;
4845: estado = 4846;
4846: estado = 4847;
4847: estado = 4848;
4848: estado = 4849;
4849: estado = 4850;
4850: estado = 4851;
4851: estado = 4852;
4852: estado = 4853;
4853: estado = 4854;
4854: estado = 4855;
4855: estado = 4856;
4856: estado = 4857;
4857: estado = 4858;
4858: estado = 4859;
4859: estado = 4860;
4860: estado = 4861;
4861: estado = 4862;
4862: estado = 4863;
4863: estado = 4864;
4864: estado = 4865;
4865: estado = 4866;
4866: estado = 4867;
4867: estado = 4868;
4868: estado = 4869;
4869: estado = 4870;
4870: estado = 4871;
4871: estado = 4872;
4872: estado = 4873;
4873: estado = 4874;
4874: estado = 4875;
4875: estado = 4876;
4876: estado = 4877;
4877: estado = 4878;
4878: estado = 4879;
4879: estado = 4880;
4880: estado = 4881;
4881: estado = 4882;
4882: estado = 4883;
4883: estado = 4884;
4884: estado = 4885;
4885: estado = 4886;
4886: estado = 4887;
4887: estado = 4888;
4888: estado = 4889;
4889: estado = 4890;
4890: estado = 4891;
4891: estado = 4892;
4892: estado = 4893;
4893: estado = 4894;
4894: estado = 4895;
4895: estado = 4896;
4896: estado = 4897;
4897: estado = 4898;
4898: estado = 4899;
4899: estado = 4900;
4900: estado = 4901;
4901: estado = 4902;
4902: estado = 4903;
4903: estado = 4904;
4904: estado = 4905;
4905: estado = 4906;
4906: estado = 4907;
4907: estado = 4908;
4908: estado = 4909;
4909: estado = 4910;
4910: estado = 4911;
4911: estado = 4912;
4912: estado = 4913;
4913: estado = 4914;
4914: estado = 4915;
4915: estado = 4916;
4916: estado = 4917;
4917: estado = 4918;
4918: estado = 4919;
4919: estado = 4920;
4920: estado = 4921;
4921: estado = 4922;
4922: estado = 4923;
4923: estado = 4924;
4924: estado = 4925;
4925: estado = 4926;
4926: estado = 4927;
4927: estado = 4928;
4928: estado = 4929;
4929: estado = 4930;
4930: estado = 4931;
4931: estado = 4932;
4932: estado = 4933;
4933: estado = 4934;
4934: estado = 4935;
4935: estado = 4936;
4936: estado = 4937;
4937: estado = 4938;
4938: estado = 4939;
4939: estado = 4940;
4940: estado = 4941;
4941: estado = 4942;
4942: estado = 4943;
4943: estado = 4944;
4944: estado = 4945;
4945: estado = 4946;
4946: estado = 4947;
4947: estado = 4948;
4948: estado = 4949;
4949: estado = 4950;
4950: estado = 4951;
4951: estado = 4952;
4952: estado = 4953;
4953: estado = 4954;
4954: estado = 4955;
4955: estado = 4956;
4956: estado = 4957;
4957: estado = 4958;
4958: estado = 4959;
4959: estado = 4960;
4960: estado = 4961;
4961: estado = 4962;
4962: estado = 4963;
4963: estado = 4964;
4964: estado = 4965;
4965: estado = 4966;
4966: estado = 4967;
4967: estado = 4968;
4968: estado = 4969;
4969: estado = 4970;
4970: estado = 4971;
4971: estado = 4972;
4972: estado = 4973;
4973: estado = 4974;
4974: estado = 4975;
4975: estado = 4976;
4976: estado = 4977;
4977: estado = 4978;
4978: estado = 4979;
4979: estado = 4980;
4980: estado = 4981;
4981: estado = 4982;
4982: estado = 4983;
4983: estado = 4984;
4984: estado = 4985;
4985: estado = 4986;
4986: estado = 4987;
4987: estado = 4988;
4988: estado = 4989;
4989: estado = 4990;
4990: estado = 4991;
4991: estado = 4992;
4992: estado = 4993;
4993: estado = 4994;
4994: estado = 4995;
4995: estado = 4996;
4996: estado = 4997;
4997: estado = 4998;
4998: estado = 4999;
4999: begin 
						estado = 5000;
						clk_out = 1;
					end
5000: estado = 5001;
5001: estado = 5002;
5002: estado = 5003;
5003: estado = 5004;
5004: estado = 5005;
5005: estado = 5006;
5006: estado = 5007;
5007: estado = 5008;
5008: estado = 5009;
5009: estado = 5010;
5010: estado = 5011;
5011: estado = 5012;
5012: estado = 5013;
5013: estado = 5014;
5014: estado = 5015;
5015: estado = 5016;
5016: estado = 5017;
5017: estado = 5018;
5018: estado = 5019;
5019: estado = 5020;
5020: estado = 5021;
5021: estado = 5022;
5022: estado = 5023;
5023: estado = 5024;
5024: estado = 5025;
5025: estado = 5026;
5026: estado = 5027;
5027: estado = 5028;
5028: estado = 5029;
5029: estado = 5030;
5030: estado = 5031;
5031: estado = 5032;
5032: estado = 5033;
5033: estado = 5034;
5034: estado = 5035;
5035: estado = 5036;
5036: estado = 5037;
5037: estado = 5038;
5038: estado = 5039;
5039: estado = 5040;
5040: estado = 5041;
5041: estado = 5042;
5042: estado = 5043;
5043: estado = 5044;
5044: estado = 5045;
5045: estado = 5046;
5046: estado = 5047;
5047: estado = 5048;
5048: estado = 5049;
5049: estado = 5050;
5050: estado = 5051;
5051: estado = 5052;
5052: estado = 5053;
5053: estado = 5054;
5054: estado = 5055;
5055: estado = 5056;
5056: estado = 5057;
5057: estado = 5058;
5058: estado = 5059;
5059: estado = 5060;
5060: estado = 5061;
5061: estado = 5062;
5062: estado = 5063;
5063: estado = 5064;
5064: estado = 5065;
5065: estado = 5066;
5066: estado = 5067;
5067: estado = 5068;
5068: estado = 5069;
5069: estado = 5070;
5070: estado = 5071;
5071: estado = 5072;
5072: estado = 5073;
5073: estado = 5074;
5074: estado = 5075;
5075: estado = 5076;
5076: estado = 5077;
5077: estado = 5078;
5078: estado = 5079;
5079: estado = 5080;
5080: estado = 5081;
5081: estado = 5082;
5082: estado = 5083;
5083: estado = 5084;
5084: estado = 5085;
5085: estado = 5086;
5086: estado = 5087;
5087: estado = 5088;
5088: estado = 5089;
5089: estado = 5090;
5090: estado = 5091;
5091: estado = 5092;
5092: estado = 5093;
5093: estado = 5094;
5094: estado = 5095;
5095: estado = 5096;
5096: estado = 5097;
5097: estado = 5098;
5098: estado = 5099;
5099: estado = 5100;
5100: estado = 5101;
5101: estado = 5102;
5102: estado = 5103;
5103: estado = 5104;
5104: estado = 5105;
5105: estado = 5106;
5106: estado = 5107;
5107: estado = 5108;
5108: estado = 5109;
5109: estado = 5110;
5110: estado = 5111;
5111: estado = 5112;
5112: estado = 5113;
5113: estado = 5114;
5114: estado = 5115;
5115: estado = 5116;
5116: estado = 5117;
5117: estado = 5118;
5118: estado = 5119;
5119: estado = 5120;
5120: estado = 5121;
5121: estado = 5122;
5122: estado = 5123;
5123: estado = 5124;
5124: estado = 5125;
5125: estado = 5126;
5126: estado = 5127;
5127: estado = 5128;
5128: estado = 5129;
5129: estado = 5130;
5130: estado = 5131;
5131: estado = 5132;
5132: estado = 5133;
5133: estado = 5134;
5134: estado = 5135;
5135: estado = 5136;
5136: estado = 5137;
5137: estado = 5138;
5138: estado = 5139;
5139: estado = 5140;
5140: estado = 5141;
5141: estado = 5142;
5142: estado = 5143;
5143: estado = 5144;
5144: estado = 5145;
5145: estado = 5146;
5146: estado = 5147;
5147: estado = 5148;
5148: estado = 5149;
5149: estado = 5150;
5150: estado = 5151;
5151: estado = 5152;
5152: estado = 5153;
5153: estado = 5154;
5154: estado = 5155;
5155: estado = 5156;
5156: estado = 5157;
5157: estado = 5158;
5158: estado = 5159;
5159: estado = 5160;
5160: estado = 5161;
5161: estado = 5162;
5162: estado = 5163;
5163: estado = 5164;
5164: estado = 5165;
5165: estado = 5166;
5166: estado = 5167;
5167: estado = 5168;
5168: estado = 5169;
5169: estado = 5170;
5170: estado = 5171;
5171: estado = 5172;
5172: estado = 5173;
5173: estado = 5174;
5174: estado = 5175;
5175: estado = 5176;
5176: estado = 5177;
5177: estado = 5178;
5178: estado = 5179;
5179: estado = 5180;
5180: estado = 5181;
5181: estado = 5182;
5182: estado = 5183;
5183: estado = 5184;
5184: estado = 5185;
5185: estado = 5186;
5186: estado = 5187;
5187: estado = 5188;
5188: estado = 5189;
5189: estado = 5190;
5190: estado = 5191;
5191: estado = 5192;
5192: estado = 5193;
5193: estado = 5194;
5194: estado = 5195;
5195: estado = 5196;
5196: estado = 5197;
5197: estado = 5198;
5198: estado = 5199;
5199: estado = 5200;
5200: estado = 5201;
5201: estado = 5202;
5202: estado = 5203;
5203: estado = 5204;
5204: estado = 5205;
5205: estado = 5206;
5206: estado = 5207;
5207: estado = 5208;
5208: estado = 5209;
5209: estado = 5210;
5210: estado = 5211;
5211: estado = 5212;
5212: estado = 5213;
5213: estado = 5214;
5214: estado = 5215;
5215: estado = 5216;
5216: estado = 5217;
5217: estado = 5218;
5218: estado = 5219;
5219: estado = 5220;
5220: estado = 5221;
5221: estado = 5222;
5222: estado = 5223;
5223: estado = 5224;
5224: estado = 5225;
5225: estado = 5226;
5226: estado = 5227;
5227: estado = 5228;
5228: estado = 5229;
5229: estado = 5230;
5230: estado = 5231;
5231: estado = 5232;
5232: estado = 5233;
5233: estado = 5234;
5234: estado = 5235;
5235: estado = 5236;
5236: estado = 5237;
5237: estado = 5238;
5238: estado = 5239;
5239: estado = 5240;
5240: estado = 5241;
5241: estado = 5242;
5242: estado = 5243;
5243: estado = 5244;
5244: estado = 5245;
5245: estado = 5246;
5246: estado = 5247;
5247: estado = 5248;
5248: estado = 5249;
5249: estado = 5250;
5250: estado = 5251;
5251: estado = 5252;
5252: estado = 5253;
5253: estado = 5254;
5254: estado = 5255;
5255: estado = 5256;
5256: estado = 5257;
5257: estado = 5258;
5258: estado = 5259;
5259: estado = 5260;
5260: estado = 5261;
5261: estado = 5262;
5262: estado = 5263;
5263: estado = 5264;
5264: estado = 5265;
5265: estado = 5266;
5266: estado = 5267;
5267: estado = 5268;
5268: estado = 5269;
5269: estado = 5270;
5270: estado = 5271;
5271: estado = 5272;
5272: estado = 5273;
5273: estado = 5274;
5274: estado = 5275;
5275: estado = 5276;
5276: estado = 5277;
5277: estado = 5278;
5278: estado = 5279;
5279: estado = 5280;
5280: estado = 5281;
5281: estado = 5282;
5282: estado = 5283;
5283: estado = 5284;
5284: estado = 5285;
5285: estado = 5286;
5286: estado = 5287;
5287: estado = 5288;
5288: estado = 5289;
5289: estado = 5290;
5290: estado = 5291;
5291: estado = 5292;
5292: estado = 5293;
5293: estado = 5294;
5294: estado = 5295;
5295: estado = 5296;
5296: estado = 5297;
5297: estado = 5298;
5298: estado = 5299;
5299: estado = 5300;
5300: estado = 5301;
5301: estado = 5302;
5302: estado = 5303;
5303: estado = 5304;
5304: estado = 5305;
5305: estado = 5306;
5306: estado = 5307;
5307: estado = 5308;
5308: estado = 5309;
5309: estado = 5310;
5310: estado = 5311;
5311: estado = 5312;
5312: estado = 5313;
5313: estado = 5314;
5314: estado = 5315;
5315: estado = 5316;
5316: estado = 5317;
5317: estado = 5318;
5318: estado = 5319;
5319: estado = 5320;
5320: estado = 5321;
5321: estado = 5322;
5322: estado = 5323;
5323: estado = 5324;
5324: estado = 5325;
5325: estado = 5326;
5326: estado = 5327;
5327: estado = 5328;
5328: estado = 5329;
5329: estado = 5330;
5330: estado = 5331;
5331: estado = 5332;
5332: estado = 5333;
5333: estado = 5334;
5334: estado = 5335;
5335: estado = 5336;
5336: estado = 5337;
5337: estado = 5338;
5338: estado = 5339;
5339: estado = 5340;
5340: estado = 5341;
5341: estado = 5342;
5342: estado = 5343;
5343: estado = 5344;
5344: estado = 5345;
5345: estado = 5346;
5346: estado = 5347;
5347: estado = 5348;
5348: estado = 5349;
5349: estado = 5350;
5350: estado = 5351;
5351: estado = 5352;
5352: estado = 5353;
5353: estado = 5354;
5354: estado = 5355;
5355: estado = 5356;
5356: estado = 5357;
5357: estado = 5358;
5358: estado = 5359;
5359: estado = 5360;
5360: estado = 5361;
5361: estado = 5362;
5362: estado = 5363;
5363: estado = 5364;
5364: estado = 5365;
5365: estado = 5366;
5366: estado = 5367;
5367: estado = 5368;
5368: estado = 5369;
5369: estado = 5370;
5370: estado = 5371;
5371: estado = 5372;
5372: estado = 5373;
5373: estado = 5374;
5374: estado = 5375;
5375: estado = 5376;
5376: estado = 5377;
5377: estado = 5378;
5378: estado = 5379;
5379: estado = 5380;
5380: estado = 5381;
5381: estado = 5382;
5382: estado = 5383;
5383: estado = 5384;
5384: estado = 5385;
5385: estado = 5386;
5386: estado = 5387;
5387: estado = 5388;
5388: estado = 5389;
5389: estado = 5390;
5390: estado = 5391;
5391: estado = 5392;
5392: estado = 5393;
5393: estado = 5394;
5394: estado = 5395;
5395: estado = 5396;
5396: estado = 5397;
5397: estado = 5398;
5398: estado = 5399;
5399: estado = 5400;
5400: estado = 5401;
5401: estado = 5402;
5402: estado = 5403;
5403: estado = 5404;
5404: estado = 5405;
5405: estado = 5406;
5406: estado = 5407;
5407: estado = 5408;
5408: estado = 5409;
5409: estado = 5410;
5410: estado = 5411;
5411: estado = 5412;
5412: estado = 5413;
5413: estado = 5414;
5414: estado = 5415;
5415: estado = 5416;
5416: estado = 5417;
5417: estado = 5418;
5418: estado = 5419;
5419: estado = 5420;
5420: estado = 5421;
5421: estado = 5422;
5422: estado = 5423;
5423: estado = 5424;
5424: estado = 5425;
5425: estado = 5426;
5426: estado = 5427;
5427: estado = 5428;
5428: estado = 5429;
5429: estado = 5430;
5430: estado = 5431;
5431: estado = 5432;
5432: estado = 5433;
5433: estado = 5434;
5434: estado = 5435;
5435: estado = 5436;
5436: estado = 5437;
5437: estado = 5438;
5438: estado = 5439;
5439: estado = 5440;
5440: estado = 5441;
5441: estado = 5442;
5442: estado = 5443;
5443: estado = 5444;
5444: estado = 5445;
5445: estado = 5446;
5446: estado = 5447;
5447: estado = 5448;
5448: estado = 5449;
5449: estado = 5450;
5450: estado = 5451;
5451: estado = 5452;
5452: estado = 5453;
5453: estado = 5454;
5454: estado = 5455;
5455: estado = 5456;
5456: estado = 5457;
5457: estado = 5458;
5458: estado = 5459;
5459: estado = 5460;
5460: estado = 5461;
5461: estado = 5462;
5462: estado = 5463;
5463: estado = 5464;
5464: estado = 5465;
5465: estado = 5466;
5466: estado = 5467;
5467: estado = 5468;
5468: estado = 5469;
5469: estado = 5470;
5470: estado = 5471;
5471: estado = 5472;
5472: estado = 5473;
5473: estado = 5474;
5474: estado = 5475;
5475: estado = 5476;
5476: estado = 5477;
5477: estado = 5478;
5478: estado = 5479;
5479: estado = 5480;
5480: estado = 5481;
5481: estado = 5482;
5482: estado = 5483;
5483: estado = 5484;
5484: estado = 5485;
5485: estado = 5486;
5486: estado = 5487;
5487: estado = 5488;
5488: estado = 5489;
5489: estado = 5490;
5490: estado = 5491;
5491: estado = 5492;
5492: estado = 5493;
5493: estado = 5494;
5494: estado = 5495;
5495: estado = 5496;
5496: estado = 5497;
5497: estado = 5498;
5498: estado = 5499;
5499: estado = 5500;
5500: estado = 5501;
5501: estado = 5502;
5502: estado = 5503;
5503: estado = 5504;
5504: estado = 5505;
5505: estado = 5506;
5506: estado = 5507;
5507: estado = 5508;
5508: estado = 5509;
5509: estado = 5510;
5510: estado = 5511;
5511: estado = 5512;
5512: estado = 5513;
5513: estado = 5514;
5514: estado = 5515;
5515: estado = 5516;
5516: estado = 5517;
5517: estado = 5518;
5518: estado = 5519;
5519: estado = 5520;
5520: estado = 5521;
5521: estado = 5522;
5522: estado = 5523;
5523: estado = 5524;
5524: estado = 5525;
5525: estado = 5526;
5526: estado = 5527;
5527: estado = 5528;
5528: estado = 5529;
5529: estado = 5530;
5530: estado = 5531;
5531: estado = 5532;
5532: estado = 5533;
5533: estado = 5534;
5534: estado = 5535;
5535: estado = 5536;
5536: estado = 5537;
5537: estado = 5538;
5538: estado = 5539;
5539: estado = 5540;
5540: estado = 5541;
5541: estado = 5542;
5542: estado = 5543;
5543: estado = 5544;
5544: estado = 5545;
5545: estado = 5546;
5546: estado = 5547;
5547: estado = 5548;
5548: estado = 5549;
5549: estado = 5550;
5550: estado = 5551;
5551: estado = 5552;
5552: estado = 5553;
5553: estado = 5554;
5554: estado = 5555;
5555: estado = 5556;
5556: estado = 5557;
5557: estado = 5558;
5558: estado = 5559;
5559: estado = 5560;
5560: estado = 5561;
5561: estado = 5562;
5562: estado = 5563;
5563: estado = 5564;
5564: estado = 5565;
5565: estado = 5566;
5566: estado = 5567;
5567: estado = 5568;
5568: estado = 5569;
5569: estado = 5570;
5570: estado = 5571;
5571: estado = 5572;
5572: estado = 5573;
5573: estado = 5574;
5574: estado = 5575;
5575: estado = 5576;
5576: estado = 5577;
5577: estado = 5578;
5578: estado = 5579;
5579: estado = 5580;
5580: estado = 5581;
5581: estado = 5582;
5582: estado = 5583;
5583: estado = 5584;
5584: estado = 5585;
5585: estado = 5586;
5586: estado = 5587;
5587: estado = 5588;
5588: estado = 5589;
5589: estado = 5590;
5590: estado = 5591;
5591: estado = 5592;
5592: estado = 5593;
5593: estado = 5594;
5594: estado = 5595;
5595: estado = 5596;
5596: estado = 5597;
5597: estado = 5598;
5598: estado = 5599;
5599: estado = 5600;
5600: estado = 5601;
5601: estado = 5602;
5602: estado = 5603;
5603: estado = 5604;
5604: estado = 5605;
5605: estado = 5606;
5606: estado = 5607;
5607: estado = 5608;
5608: estado = 5609;
5609: estado = 5610;
5610: estado = 5611;
5611: estado = 5612;
5612: estado = 5613;
5613: estado = 5614;
5614: estado = 5615;
5615: estado = 5616;
5616: estado = 5617;
5617: estado = 5618;
5618: estado = 5619;
5619: estado = 5620;
5620: estado = 5621;
5621: estado = 5622;
5622: estado = 5623;
5623: estado = 5624;
5624: estado = 5625;
5625: estado = 5626;
5626: estado = 5627;
5627: estado = 5628;
5628: estado = 5629;
5629: estado = 5630;
5630: estado = 5631;
5631: estado = 5632;
5632: estado = 5633;
5633: estado = 5634;
5634: estado = 5635;
5635: estado = 5636;
5636: estado = 5637;
5637: estado = 5638;
5638: estado = 5639;
5639: estado = 5640;
5640: estado = 5641;
5641: estado = 5642;
5642: estado = 5643;
5643: estado = 5644;
5644: estado = 5645;
5645: estado = 5646;
5646: estado = 5647;
5647: estado = 5648;
5648: estado = 5649;
5649: estado = 5650;
5650: estado = 5651;
5651: estado = 5652;
5652: estado = 5653;
5653: estado = 5654;
5654: estado = 5655;
5655: estado = 5656;
5656: estado = 5657;
5657: estado = 5658;
5658: estado = 5659;
5659: estado = 5660;
5660: estado = 5661;
5661: estado = 5662;
5662: estado = 5663;
5663: estado = 5664;
5664: estado = 5665;
5665: estado = 5666;
5666: estado = 5667;
5667: estado = 5668;
5668: estado = 5669;
5669: estado = 5670;
5670: estado = 5671;
5671: estado = 5672;
5672: estado = 5673;
5673: estado = 5674;
5674: estado = 5675;
5675: estado = 5676;
5676: estado = 5677;
5677: estado = 5678;
5678: estado = 5679;
5679: estado = 5680;
5680: estado = 5681;
5681: estado = 5682;
5682: estado = 5683;
5683: estado = 5684;
5684: estado = 5685;
5685: estado = 5686;
5686: estado = 5687;
5687: estado = 5688;
5688: estado = 5689;
5689: estado = 5690;
5690: estado = 5691;
5691: estado = 5692;
5692: estado = 5693;
5693: estado = 5694;
5694: estado = 5695;
5695: estado = 5696;
5696: estado = 5697;
5697: estado = 5698;
5698: estado = 5699;
5699: estado = 5700;
5700: estado = 5701;
5701: estado = 5702;
5702: estado = 5703;
5703: estado = 5704;
5704: estado = 5705;
5705: estado = 5706;
5706: estado = 5707;
5707: estado = 5708;
5708: estado = 5709;
5709: estado = 5710;
5710: estado = 5711;
5711: estado = 5712;
5712: estado = 5713;
5713: estado = 5714;
5714: estado = 5715;
5715: estado = 5716;
5716: estado = 5717;
5717: estado = 5718;
5718: estado = 5719;
5719: estado = 5720;
5720: estado = 5721;
5721: estado = 5722;
5722: estado = 5723;
5723: estado = 5724;
5724: estado = 5725;
5725: estado = 5726;
5726: estado = 5727;
5727: estado = 5728;
5728: estado = 5729;
5729: estado = 5730;
5730: estado = 5731;
5731: estado = 5732;
5732: estado = 5733;
5733: estado = 5734;
5734: estado = 5735;
5735: estado = 5736;
5736: estado = 5737;
5737: estado = 5738;
5738: estado = 5739;
5739: estado = 5740;
5740: estado = 5741;
5741: estado = 5742;
5742: estado = 5743;
5743: estado = 5744;
5744: estado = 5745;
5745: estado = 5746;
5746: estado = 5747;
5747: estado = 5748;
5748: estado = 5749;
5749: estado = 5750;
5750: estado = 5751;
5751: estado = 5752;
5752: estado = 5753;
5753: estado = 5754;
5754: estado = 5755;
5755: estado = 5756;
5756: estado = 5757;
5757: estado = 5758;
5758: estado = 5759;
5759: estado = 5760;
5760: estado = 5761;
5761: estado = 5762;
5762: estado = 5763;
5763: estado = 5764;
5764: estado = 5765;
5765: estado = 5766;
5766: estado = 5767;
5767: estado = 5768;
5768: estado = 5769;
5769: estado = 5770;
5770: estado = 5771;
5771: estado = 5772;
5772: estado = 5773;
5773: estado = 5774;
5774: estado = 5775;
5775: estado = 5776;
5776: estado = 5777;
5777: estado = 5778;
5778: estado = 5779;
5779: estado = 5780;
5780: estado = 5781;
5781: estado = 5782;
5782: estado = 5783;
5783: estado = 5784;
5784: estado = 5785;
5785: estado = 5786;
5786: estado = 5787;
5787: estado = 5788;
5788: estado = 5789;
5789: estado = 5790;
5790: estado = 5791;
5791: estado = 5792;
5792: estado = 5793;
5793: estado = 5794;
5794: estado = 5795;
5795: estado = 5796;
5796: estado = 5797;
5797: estado = 5798;
5798: estado = 5799;
5799: estado = 5800;
5800: estado = 5801;
5801: estado = 5802;
5802: estado = 5803;
5803: estado = 5804;
5804: estado = 5805;
5805: estado = 5806;
5806: estado = 5807;
5807: estado = 5808;
5808: estado = 5809;
5809: estado = 5810;
5810: estado = 5811;
5811: estado = 5812;
5812: estado = 5813;
5813: estado = 5814;
5814: estado = 5815;
5815: estado = 5816;
5816: estado = 5817;
5817: estado = 5818;
5818: estado = 5819;
5819: estado = 5820;
5820: estado = 5821;
5821: estado = 5822;
5822: estado = 5823;
5823: estado = 5824;
5824: estado = 5825;
5825: estado = 5826;
5826: estado = 5827;
5827: estado = 5828;
5828: estado = 5829;
5829: estado = 5830;
5830: estado = 5831;
5831: estado = 5832;
5832: estado = 5833;
5833: estado = 5834;
5834: estado = 5835;
5835: estado = 5836;
5836: estado = 5837;
5837: estado = 5838;
5838: estado = 5839;
5839: estado = 5840;
5840: estado = 5841;
5841: estado = 5842;
5842: estado = 5843;
5843: estado = 5844;
5844: estado = 5845;
5845: estado = 5846;
5846: estado = 5847;
5847: estado = 5848;
5848: estado = 5849;
5849: estado = 5850;
5850: estado = 5851;
5851: estado = 5852;
5852: estado = 5853;
5853: estado = 5854;
5854: estado = 5855;
5855: estado = 5856;
5856: estado = 5857;
5857: estado = 5858;
5858: estado = 5859;
5859: estado = 5860;
5860: estado = 5861;
5861: estado = 5862;
5862: estado = 5863;
5863: estado = 5864;
5864: estado = 5865;
5865: estado = 5866;
5866: estado = 5867;
5867: estado = 5868;
5868: estado = 5869;
5869: estado = 5870;
5870: estado = 5871;
5871: estado = 5872;
5872: estado = 5873;
5873: estado = 5874;
5874: estado = 5875;
5875: estado = 5876;
5876: estado = 5877;
5877: estado = 5878;
5878: estado = 5879;
5879: estado = 5880;
5880: estado = 5881;
5881: estado = 5882;
5882: estado = 5883;
5883: estado = 5884;
5884: estado = 5885;
5885: estado = 5886;
5886: estado = 5887;
5887: estado = 5888;
5888: estado = 5889;
5889: estado = 5890;
5890: estado = 5891;
5891: estado = 5892;
5892: estado = 5893;
5893: estado = 5894;
5894: estado = 5895;
5895: estado = 5896;
5896: estado = 5897;
5897: estado = 5898;
5898: estado = 5899;
5899: estado = 5900;
5900: estado = 5901;
5901: estado = 5902;
5902: estado = 5903;
5903: estado = 5904;
5904: estado = 5905;
5905: estado = 5906;
5906: estado = 5907;
5907: estado = 5908;
5908: estado = 5909;
5909: estado = 5910;
5910: estado = 5911;
5911: estado = 5912;
5912: estado = 5913;
5913: estado = 5914;
5914: estado = 5915;
5915: estado = 5916;
5916: estado = 5917;
5917: estado = 5918;
5918: estado = 5919;
5919: estado = 5920;
5920: estado = 5921;
5921: estado = 5922;
5922: estado = 5923;
5923: estado = 5924;
5924: estado = 5925;
5925: estado = 5926;
5926: estado = 5927;
5927: estado = 5928;
5928: estado = 5929;
5929: estado = 5930;
5930: estado = 5931;
5931: estado = 5932;
5932: estado = 5933;
5933: estado = 5934;
5934: estado = 5935;
5935: estado = 5936;
5936: estado = 5937;
5937: estado = 5938;
5938: estado = 5939;
5939: estado = 5940;
5940: estado = 5941;
5941: estado = 5942;
5942: estado = 5943;
5943: estado = 5944;
5944: estado = 5945;
5945: estado = 5946;
5946: estado = 5947;
5947: estado = 5948;
5948: estado = 5949;
5949: estado = 5950;
5950: estado = 5951;
5951: estado = 5952;
5952: estado = 5953;
5953: estado = 5954;
5954: estado = 5955;
5955: estado = 5956;
5956: estado = 5957;
5957: estado = 5958;
5958: estado = 5959;
5959: estado = 5960;
5960: estado = 5961;
5961: estado = 5962;
5962: estado = 5963;
5963: estado = 5964;
5964: estado = 5965;
5965: estado = 5966;
5966: estado = 5967;
5967: estado = 5968;
5968: estado = 5969;
5969: estado = 5970;
5970: estado = 5971;
5971: estado = 5972;
5972: estado = 5973;
5973: estado = 5974;
5974: estado = 5975;
5975: estado = 5976;
5976: estado = 5977;
5977: estado = 5978;
5978: estado = 5979;
5979: estado = 5980;
5980: estado = 5981;
5981: estado = 5982;
5982: estado = 5983;
5983: estado = 5984;
5984: estado = 5985;
5985: estado = 5986;
5986: estado = 5987;
5987: estado = 5988;
5988: estado = 5989;
5989: estado = 5990;
5990: estado = 5991;
5991: estado = 5992;
5992: estado = 5993;
5993: estado = 5994;
5994: estado = 5995;
5995: estado = 5996;
5996: estado = 5997;
5997: estado = 5998;
5998: estado = 5999;
5999: estado = 6000;
6000: estado = 6001;
6001: estado = 6002;
6002: estado = 6003;
6003: estado = 6004;
6004: estado = 6005;
6005: estado = 6006;
6006: estado = 6007;
6007: estado = 6008;
6008: estado = 6009;
6009: estado = 6010;
6010: estado = 6011;
6011: estado = 6012;
6012: estado = 6013;
6013: estado = 6014;
6014: estado = 6015;
6015: estado = 6016;
6016: estado = 6017;
6017: estado = 6018;
6018: estado = 6019;
6019: estado = 6020;
6020: estado = 6021;
6021: estado = 6022;
6022: estado = 6023;
6023: estado = 6024;
6024: estado = 6025;
6025: estado = 6026;
6026: estado = 6027;
6027: estado = 6028;
6028: estado = 6029;
6029: estado = 6030;
6030: estado = 6031;
6031: estado = 6032;
6032: estado = 6033;
6033: estado = 6034;
6034: estado = 6035;
6035: estado = 6036;
6036: estado = 6037;
6037: estado = 6038;
6038: estado = 6039;
6039: estado = 6040;
6040: estado = 6041;
6041: estado = 6042;
6042: estado = 6043;
6043: estado = 6044;
6044: estado = 6045;
6045: estado = 6046;
6046: estado = 6047;
6047: estado = 6048;
6048: estado = 6049;
6049: estado = 6050;
6050: estado = 6051;
6051: estado = 6052;
6052: estado = 6053;
6053: estado = 6054;
6054: estado = 6055;
6055: estado = 6056;
6056: estado = 6057;
6057: estado = 6058;
6058: estado = 6059;
6059: estado = 6060;
6060: estado = 6061;
6061: estado = 6062;
6062: estado = 6063;
6063: estado = 6064;
6064: estado = 6065;
6065: estado = 6066;
6066: estado = 6067;
6067: estado = 6068;
6068: estado = 6069;
6069: estado = 6070;
6070: estado = 6071;
6071: estado = 6072;
6072: estado = 6073;
6073: estado = 6074;
6074: estado = 6075;
6075: estado = 6076;
6076: estado = 6077;
6077: estado = 6078;
6078: estado = 6079;
6079: estado = 6080;
6080: estado = 6081;
6081: estado = 6082;
6082: estado = 6083;
6083: estado = 6084;
6084: estado = 6085;
6085: estado = 6086;
6086: estado = 6087;
6087: estado = 6088;
6088: estado = 6089;
6089: estado = 6090;
6090: estado = 6091;
6091: estado = 6092;
6092: estado = 6093;
6093: estado = 6094;
6094: estado = 6095;
6095: estado = 6096;
6096: estado = 6097;
6097: estado = 6098;
6098: estado = 6099;
6099: estado = 6100;
6100: estado = 6101;
6101: estado = 6102;
6102: estado = 6103;
6103: estado = 6104;
6104: estado = 6105;
6105: estado = 6106;
6106: estado = 6107;
6107: estado = 6108;
6108: estado = 6109;
6109: estado = 6110;
6110: estado = 6111;
6111: estado = 6112;
6112: estado = 6113;
6113: estado = 6114;
6114: estado = 6115;
6115: estado = 6116;
6116: estado = 6117;
6117: estado = 6118;
6118: estado = 6119;
6119: estado = 6120;
6120: estado = 6121;
6121: estado = 6122;
6122: estado = 6123;
6123: estado = 6124;
6124: estado = 6125;
6125: estado = 6126;
6126: estado = 6127;
6127: estado = 6128;
6128: estado = 6129;
6129: estado = 6130;
6130: estado = 6131;
6131: estado = 6132;
6132: estado = 6133;
6133: estado = 6134;
6134: estado = 6135;
6135: estado = 6136;
6136: estado = 6137;
6137: estado = 6138;
6138: estado = 6139;
6139: estado = 6140;
6140: estado = 6141;
6141: estado = 6142;
6142: estado = 6143;
6143: estado = 6144;
6144: estado = 6145;
6145: estado = 6146;
6146: estado = 6147;
6147: estado = 6148;
6148: estado = 6149;
6149: estado = 6150;
6150: estado = 6151;
6151: estado = 6152;
6152: estado = 6153;
6153: estado = 6154;
6154: estado = 6155;
6155: estado = 6156;
6156: estado = 6157;
6157: estado = 6158;
6158: estado = 6159;
6159: estado = 6160;
6160: estado = 6161;
6161: estado = 6162;
6162: estado = 6163;
6163: estado = 6164;
6164: estado = 6165;
6165: estado = 6166;
6166: estado = 6167;
6167: estado = 6168;
6168: estado = 6169;
6169: estado = 6170;
6170: estado = 6171;
6171: estado = 6172;
6172: estado = 6173;
6173: estado = 6174;
6174: estado = 6175;
6175: estado = 6176;
6176: estado = 6177;
6177: estado = 6178;
6178: estado = 6179;
6179: estado = 6180;
6180: estado = 6181;
6181: estado = 6182;
6182: estado = 6183;
6183: estado = 6184;
6184: estado = 6185;
6185: estado = 6186;
6186: estado = 6187;
6187: estado = 6188;
6188: estado = 6189;
6189: estado = 6190;
6190: estado = 6191;
6191: estado = 6192;
6192: estado = 6193;
6193: estado = 6194;
6194: estado = 6195;
6195: estado = 6196;
6196: estado = 6197;
6197: estado = 6198;
6198: estado = 6199;
6199: estado = 6200;
6200: estado = 6201;
6201: estado = 6202;
6202: estado = 6203;
6203: estado = 6204;
6204: estado = 6205;
6205: estado = 6206;
6206: estado = 6207;
6207: estado = 6208;
6208: estado = 6209;
6209: estado = 6210;
6210: estado = 6211;
6211: estado = 6212;
6212: estado = 6213;
6213: estado = 6214;
6214: estado = 6215;
6215: estado = 6216;
6216: estado = 6217;
6217: estado = 6218;
6218: estado = 6219;
6219: estado = 6220;
6220: estado = 6221;
6221: estado = 6222;
6222: estado = 6223;
6223: estado = 6224;
6224: estado = 6225;
6225: estado = 6226;
6226: estado = 6227;
6227: estado = 6228;
6228: estado = 6229;
6229: estado = 6230;
6230: estado = 6231;
6231: estado = 6232;
6232: estado = 6233;
6233: estado = 6234;
6234: estado = 6235;
6235: estado = 6236;
6236: estado = 6237;
6237: estado = 6238;
6238: estado = 6239;
6239: estado = 6240;
6240: estado = 6241;
6241: estado = 6242;
6242: estado = 6243;
6243: estado = 6244;
6244: estado = 6245;
6245: estado = 6246;
6246: estado = 6247;
6247: estado = 6248;
6248: estado = 6249;
6249: estado = 6250;
6250: estado = 6251;
6251: estado = 6252;
6252: estado = 6253;
6253: estado = 6254;
6254: estado = 6255;
6255: estado = 6256;
6256: estado = 6257;
6257: estado = 6258;
6258: estado = 6259;
6259: estado = 6260;
6260: estado = 6261;
6261: estado = 6262;
6262: estado = 6263;
6263: estado = 6264;
6264: estado = 6265;
6265: estado = 6266;
6266: estado = 6267;
6267: estado = 6268;
6268: estado = 6269;
6269: estado = 6270;
6270: estado = 6271;
6271: estado = 6272;
6272: estado = 6273;
6273: estado = 6274;
6274: estado = 6275;
6275: estado = 6276;
6276: estado = 6277;
6277: estado = 6278;
6278: estado = 6279;
6279: estado = 6280;
6280: estado = 6281;
6281: estado = 6282;
6282: estado = 6283;
6283: estado = 6284;
6284: estado = 6285;
6285: estado = 6286;
6286: estado = 6287;
6287: estado = 6288;
6288: estado = 6289;
6289: estado = 6290;
6290: estado = 6291;
6291: estado = 6292;
6292: estado = 6293;
6293: estado = 6294;
6294: estado = 6295;
6295: estado = 6296;
6296: estado = 6297;
6297: estado = 6298;
6298: estado = 6299;
6299: estado = 6300;
6300: estado = 6301;
6301: estado = 6302;
6302: estado = 6303;
6303: estado = 6304;
6304: estado = 6305;
6305: estado = 6306;
6306: estado = 6307;
6307: estado = 6308;
6308: estado = 6309;
6309: estado = 6310;
6310: estado = 6311;
6311: estado = 6312;
6312: estado = 6313;
6313: estado = 6314;
6314: estado = 6315;
6315: estado = 6316;
6316: estado = 6317;
6317: estado = 6318;
6318: estado = 6319;
6319: estado = 6320;
6320: estado = 6321;
6321: estado = 6322;
6322: estado = 6323;
6323: estado = 6324;
6324: estado = 6325;
6325: estado = 6326;
6326: estado = 6327;
6327: estado = 6328;
6328: estado = 6329;
6329: estado = 6330;
6330: estado = 6331;
6331: estado = 6332;
6332: estado = 6333;
6333: estado = 6334;
6334: estado = 6335;
6335: estado = 6336;
6336: estado = 6337;
6337: estado = 6338;
6338: estado = 6339;
6339: estado = 6340;
6340: estado = 6341;
6341: estado = 6342;
6342: estado = 6343;
6343: estado = 6344;
6344: estado = 6345;
6345: estado = 6346;
6346: estado = 6347;
6347: estado = 6348;
6348: estado = 6349;
6349: estado = 6350;
6350: estado = 6351;
6351: estado = 6352;
6352: estado = 6353;
6353: estado = 6354;
6354: estado = 6355;
6355: estado = 6356;
6356: estado = 6357;
6357: estado = 6358;
6358: estado = 6359;
6359: estado = 6360;
6360: estado = 6361;
6361: estado = 6362;
6362: estado = 6363;
6363: estado = 6364;
6364: estado = 6365;
6365: estado = 6366;
6366: estado = 6367;
6367: estado = 6368;
6368: estado = 6369;
6369: estado = 6370;
6370: estado = 6371;
6371: estado = 6372;
6372: estado = 6373;
6373: estado = 6374;
6374: estado = 6375;
6375: estado = 6376;
6376: estado = 6377;
6377: estado = 6378;
6378: estado = 6379;
6379: estado = 6380;
6380: estado = 6381;
6381: estado = 6382;
6382: estado = 6383;
6383: estado = 6384;
6384: estado = 6385;
6385: estado = 6386;
6386: estado = 6387;
6387: estado = 6388;
6388: estado = 6389;
6389: estado = 6390;
6390: estado = 6391;
6391: estado = 6392;
6392: estado = 6393;
6393: estado = 6394;
6394: estado = 6395;
6395: estado = 6396;
6396: estado = 6397;
6397: estado = 6398;
6398: estado = 6399;
6399: estado = 6400;
6400: estado = 6401;
6401: estado = 6402;
6402: estado = 6403;
6403: estado = 6404;
6404: estado = 6405;
6405: estado = 6406;
6406: estado = 6407;
6407: estado = 6408;
6408: estado = 6409;
6409: estado = 6410;
6410: estado = 6411;
6411: estado = 6412;
6412: estado = 6413;
6413: estado = 6414;
6414: estado = 6415;
6415: estado = 6416;
6416: estado = 6417;
6417: estado = 6418;
6418: estado = 6419;
6419: estado = 6420;
6420: estado = 6421;
6421: estado = 6422;
6422: estado = 6423;
6423: estado = 6424;
6424: estado = 6425;
6425: estado = 6426;
6426: estado = 6427;
6427: estado = 6428;
6428: estado = 6429;
6429: estado = 6430;
6430: estado = 6431;
6431: estado = 6432;
6432: estado = 6433;
6433: estado = 6434;
6434: estado = 6435;
6435: estado = 6436;
6436: estado = 6437;
6437: estado = 6438;
6438: estado = 6439;
6439: estado = 6440;
6440: estado = 6441;
6441: estado = 6442;
6442: estado = 6443;
6443: estado = 6444;
6444: estado = 6445;
6445: estado = 6446;
6446: estado = 6447;
6447: estado = 6448;
6448: estado = 6449;
6449: estado = 6450;
6450: estado = 6451;
6451: estado = 6452;
6452: estado = 6453;
6453: estado = 6454;
6454: estado = 6455;
6455: estado = 6456;
6456: estado = 6457;
6457: estado = 6458;
6458: estado = 6459;
6459: estado = 6460;
6460: estado = 6461;
6461: estado = 6462;
6462: estado = 6463;
6463: estado = 6464;
6464: estado = 6465;
6465: estado = 6466;
6466: estado = 6467;
6467: estado = 6468;
6468: estado = 6469;
6469: estado = 6470;
6470: estado = 6471;
6471: estado = 6472;
6472: estado = 6473;
6473: estado = 6474;
6474: estado = 6475;
6475: estado = 6476;
6476: estado = 6477;
6477: estado = 6478;
6478: estado = 6479;
6479: estado = 6480;
6480: estado = 6481;
6481: estado = 6482;
6482: estado = 6483;
6483: estado = 6484;
6484: estado = 6485;
6485: estado = 6486;
6486: estado = 6487;
6487: estado = 6488;
6488: estado = 6489;
6489: estado = 6490;
6490: estado = 6491;
6491: estado = 6492;
6492: estado = 6493;
6493: estado = 6494;
6494: estado = 6495;
6495: estado = 6496;
6496: estado = 6497;
6497: estado = 6498;
6498: estado = 6499;
6499: estado = 6500;
6500: estado = 6501;
6501: estado = 6502;
6502: estado = 6503;
6503: estado = 6504;
6504: estado = 6505;
6505: estado = 6506;
6506: estado = 6507;
6507: estado = 6508;
6508: estado = 6509;
6509: estado = 6510;
6510: estado = 6511;
6511: estado = 6512;
6512: estado = 6513;
6513: estado = 6514;
6514: estado = 6515;
6515: estado = 6516;
6516: estado = 6517;
6517: estado = 6518;
6518: estado = 6519;
6519: estado = 6520;
6520: estado = 6521;
6521: estado = 6522;
6522: estado = 6523;
6523: estado = 6524;
6524: estado = 6525;
6525: estado = 6526;
6526: estado = 6527;
6527: estado = 6528;
6528: estado = 6529;
6529: estado = 6530;
6530: estado = 6531;
6531: estado = 6532;
6532: estado = 6533;
6533: estado = 6534;
6534: estado = 6535;
6535: estado = 6536;
6536: estado = 6537;
6537: estado = 6538;
6538: estado = 6539;
6539: estado = 6540;
6540: estado = 6541;
6541: estado = 6542;
6542: estado = 6543;
6543: estado = 6544;
6544: estado = 6545;
6545: estado = 6546;
6546: estado = 6547;
6547: estado = 6548;
6548: estado = 6549;
6549: estado = 6550;
6550: estado = 6551;
6551: estado = 6552;
6552: estado = 6553;
6553: estado = 6554;
6554: estado = 6555;
6555: estado = 6556;
6556: estado = 6557;
6557: estado = 6558;
6558: estado = 6559;
6559: estado = 6560;
6560: estado = 6561;
6561: estado = 6562;
6562: estado = 6563;
6563: estado = 6564;
6564: estado = 6565;
6565: estado = 6566;
6566: estado = 6567;
6567: estado = 6568;
6568: estado = 6569;
6569: estado = 6570;
6570: estado = 6571;
6571: estado = 6572;
6572: estado = 6573;
6573: estado = 6574;
6574: estado = 6575;
6575: estado = 6576;
6576: estado = 6577;
6577: estado = 6578;
6578: estado = 6579;
6579: estado = 6580;
6580: estado = 6581;
6581: estado = 6582;
6582: estado = 6583;
6583: estado = 6584;
6584: estado = 6585;
6585: estado = 6586;
6586: estado = 6587;
6587: estado = 6588;
6588: estado = 6589;
6589: estado = 6590;
6590: estado = 6591;
6591: estado = 6592;
6592: estado = 6593;
6593: estado = 6594;
6594: estado = 6595;
6595: estado = 6596;
6596: estado = 6597;
6597: estado = 6598;
6598: estado = 6599;
6599: estado = 6600;
6600: estado = 6601;
6601: estado = 6602;
6602: estado = 6603;
6603: estado = 6604;
6604: estado = 6605;
6605: estado = 6606;
6606: estado = 6607;
6607: estado = 6608;
6608: estado = 6609;
6609: estado = 6610;
6610: estado = 6611;
6611: estado = 6612;
6612: estado = 6613;
6613: estado = 6614;
6614: estado = 6615;
6615: estado = 6616;
6616: estado = 6617;
6617: estado = 6618;
6618: estado = 6619;
6619: estado = 6620;
6620: estado = 6621;
6621: estado = 6622;
6622: estado = 6623;
6623: estado = 6624;
6624: estado = 6625;
6625: estado = 6626;
6626: estado = 6627;
6627: estado = 6628;
6628: estado = 6629;
6629: estado = 6630;
6630: estado = 6631;
6631: estado = 6632;
6632: estado = 6633;
6633: estado = 6634;
6634: estado = 6635;
6635: estado = 6636;
6636: estado = 6637;
6637: estado = 6638;
6638: estado = 6639;
6639: estado = 6640;
6640: estado = 6641;
6641: estado = 6642;
6642: estado = 6643;
6643: estado = 6644;
6644: estado = 6645;
6645: estado = 6646;
6646: estado = 6647;
6647: estado = 6648;
6648: estado = 6649;
6649: estado = 6650;
6650: estado = 6651;
6651: estado = 6652;
6652: estado = 6653;
6653: estado = 6654;
6654: estado = 6655;
6655: estado = 6656;
6656: estado = 6657;
6657: estado = 6658;
6658: estado = 6659;
6659: estado = 6660;
6660: estado = 6661;
6661: estado = 6662;
6662: estado = 6663;
6663: estado = 6664;
6664: estado = 6665;
6665: estado = 6666;
6666: estado = 6667;
6667: estado = 6668;
6668: estado = 6669;
6669: estado = 6670;
6670: estado = 6671;
6671: estado = 6672;
6672: estado = 6673;
6673: estado = 6674;
6674: estado = 6675;
6675: estado = 6676;
6676: estado = 6677;
6677: estado = 6678;
6678: estado = 6679;
6679: estado = 6680;
6680: estado = 6681;
6681: estado = 6682;
6682: estado = 6683;
6683: estado = 6684;
6684: estado = 6685;
6685: estado = 6686;
6686: estado = 6687;
6687: estado = 6688;
6688: estado = 6689;
6689: estado = 6690;
6690: estado = 6691;
6691: estado = 6692;
6692: estado = 6693;
6693: estado = 6694;
6694: estado = 6695;
6695: estado = 6696;
6696: estado = 6697;
6697: estado = 6698;
6698: estado = 6699;
6699: estado = 6700;
6700: estado = 6701;
6701: estado = 6702;
6702: estado = 6703;
6703: estado = 6704;
6704: estado = 6705;
6705: estado = 6706;
6706: estado = 6707;
6707: estado = 6708;
6708: estado = 6709;
6709: estado = 6710;
6710: estado = 6711;
6711: estado = 6712;
6712: estado = 6713;
6713: estado = 6714;
6714: estado = 6715;
6715: estado = 6716;
6716: estado = 6717;
6717: estado = 6718;
6718: estado = 6719;
6719: estado = 6720;
6720: estado = 6721;
6721: estado = 6722;
6722: estado = 6723;
6723: estado = 6724;
6724: estado = 6725;
6725: estado = 6726;
6726: estado = 6727;
6727: estado = 6728;
6728: estado = 6729;
6729: estado = 6730;
6730: estado = 6731;
6731: estado = 6732;
6732: estado = 6733;
6733: estado = 6734;
6734: estado = 6735;
6735: estado = 6736;
6736: estado = 6737;
6737: estado = 6738;
6738: estado = 6739;
6739: estado = 6740;
6740: estado = 6741;
6741: estado = 6742;
6742: estado = 6743;
6743: estado = 6744;
6744: estado = 6745;
6745: estado = 6746;
6746: estado = 6747;
6747: estado = 6748;
6748: estado = 6749;
6749: estado = 6750;
6750: estado = 6751;
6751: estado = 6752;
6752: estado = 6753;
6753: estado = 6754;
6754: estado = 6755;
6755: estado = 6756;
6756: estado = 6757;
6757: estado = 6758;
6758: estado = 6759;
6759: estado = 6760;
6760: estado = 6761;
6761: estado = 6762;
6762: estado = 6763;
6763: estado = 6764;
6764: estado = 6765;
6765: estado = 6766;
6766: estado = 6767;
6767: estado = 6768;
6768: estado = 6769;
6769: estado = 6770;
6770: estado = 6771;
6771: estado = 6772;
6772: estado = 6773;
6773: estado = 6774;
6774: estado = 6775;
6775: estado = 6776;
6776: estado = 6777;
6777: estado = 6778;
6778: estado = 6779;
6779: estado = 6780;
6780: estado = 6781;
6781: estado = 6782;
6782: estado = 6783;
6783: estado = 6784;
6784: estado = 6785;
6785: estado = 6786;
6786: estado = 6787;
6787: estado = 6788;
6788: estado = 6789;
6789: estado = 6790;
6790: estado = 6791;
6791: estado = 6792;
6792: estado = 6793;
6793: estado = 6794;
6794: estado = 6795;
6795: estado = 6796;
6796: estado = 6797;
6797: estado = 6798;
6798: estado = 6799;
6799: estado = 6800;
6800: estado = 6801;
6801: estado = 6802;
6802: estado = 6803;
6803: estado = 6804;
6804: estado = 6805;
6805: estado = 6806;
6806: estado = 6807;
6807: estado = 6808;
6808: estado = 6809;
6809: estado = 6810;
6810: estado = 6811;
6811: estado = 6812;
6812: estado = 6813;
6813: estado = 6814;
6814: estado = 6815;
6815: estado = 6816;
6816: estado = 6817;
6817: estado = 6818;
6818: estado = 6819;
6819: estado = 6820;
6820: estado = 6821;
6821: estado = 6822;
6822: estado = 6823;
6823: estado = 6824;
6824: estado = 6825;
6825: estado = 6826;
6826: estado = 6827;
6827: estado = 6828;
6828: estado = 6829;
6829: estado = 6830;
6830: estado = 6831;
6831: estado = 6832;
6832: estado = 6833;
6833: estado = 6834;
6834: estado = 6835;
6835: estado = 6836;
6836: estado = 6837;
6837: estado = 6838;
6838: estado = 6839;
6839: estado = 6840;
6840: estado = 6841;
6841: estado = 6842;
6842: estado = 6843;
6843: estado = 6844;
6844: estado = 6845;
6845: estado = 6846;
6846: estado = 6847;
6847: estado = 6848;
6848: estado = 6849;
6849: estado = 6850;
6850: estado = 6851;
6851: estado = 6852;
6852: estado = 6853;
6853: estado = 6854;
6854: estado = 6855;
6855: estado = 6856;
6856: estado = 6857;
6857: estado = 6858;
6858: estado = 6859;
6859: estado = 6860;
6860: estado = 6861;
6861: estado = 6862;
6862: estado = 6863;
6863: estado = 6864;
6864: estado = 6865;
6865: estado = 6866;
6866: estado = 6867;
6867: estado = 6868;
6868: estado = 6869;
6869: estado = 6870;
6870: estado = 6871;
6871: estado = 6872;
6872: estado = 6873;
6873: estado = 6874;
6874: estado = 6875;
6875: estado = 6876;
6876: estado = 6877;
6877: estado = 6878;
6878: estado = 6879;
6879: estado = 6880;
6880: estado = 6881;
6881: estado = 6882;
6882: estado = 6883;
6883: estado = 6884;
6884: estado = 6885;
6885: estado = 6886;
6886: estado = 6887;
6887: estado = 6888;
6888: estado = 6889;
6889: estado = 6890;
6890: estado = 6891;
6891: estado = 6892;
6892: estado = 6893;
6893: estado = 6894;
6894: estado = 6895;
6895: estado = 6896;
6896: estado = 6897;
6897: estado = 6898;
6898: estado = 6899;
6899: estado = 6900;
6900: estado = 6901;
6901: estado = 6902;
6902: estado = 6903;
6903: estado = 6904;
6904: estado = 6905;
6905: estado = 6906;
6906: estado = 6907;
6907: estado = 6908;
6908: estado = 6909;
6909: estado = 6910;
6910: estado = 6911;
6911: estado = 6912;
6912: estado = 6913;
6913: estado = 6914;
6914: estado = 6915;
6915: estado = 6916;
6916: estado = 6917;
6917: estado = 6918;
6918: estado = 6919;
6919: estado = 6920;
6920: estado = 6921;
6921: estado = 6922;
6922: estado = 6923;
6923: estado = 6924;
6924: estado = 6925;
6925: estado = 6926;
6926: estado = 6927;
6927: estado = 6928;
6928: estado = 6929;
6929: estado = 6930;
6930: estado = 6931;
6931: estado = 6932;
6932: estado = 6933;
6933: estado = 6934;
6934: estado = 6935;
6935: estado = 6936;
6936: estado = 6937;
6937: estado = 6938;
6938: estado = 6939;
6939: estado = 6940;
6940: estado = 6941;
6941: estado = 6942;
6942: estado = 6943;
6943: estado = 6944;
6944: estado = 6945;
6945: estado = 6946;
6946: estado = 6947;
6947: estado = 6948;
6948: estado = 6949;
6949: estado = 6950;
6950: estado = 6951;
6951: estado = 6952;
6952: estado = 6953;
6953: estado = 6954;
6954: estado = 6955;
6955: estado = 6956;
6956: estado = 6957;
6957: estado = 6958;
6958: estado = 6959;
6959: estado = 6960;
6960: estado = 6961;
6961: estado = 6962;
6962: estado = 6963;
6963: estado = 6964;
6964: estado = 6965;
6965: estado = 6966;
6966: estado = 6967;
6967: estado = 6968;
6968: estado = 6969;
6969: estado = 6970;
6970: estado = 6971;
6971: estado = 6972;
6972: estado = 6973;
6973: estado = 6974;
6974: estado = 6975;
6975: estado = 6976;
6976: estado = 6977;
6977: estado = 6978;
6978: estado = 6979;
6979: estado = 6980;
6980: estado = 6981;
6981: estado = 6982;
6982: estado = 6983;
6983: estado = 6984;
6984: estado = 6985;
6985: estado = 6986;
6986: estado = 6987;
6987: estado = 6988;
6988: estado = 6989;
6989: estado = 6990;
6990: estado = 6991;
6991: estado = 6992;
6992: estado = 6993;
6993: estado = 6994;
6994: estado = 6995;
6995: estado = 6996;
6996: estado = 6997;
6997: estado = 6998;
6998: estado = 6999;
6999: estado = 7000;
7000: estado = 7001;
7001: estado = 7002;
7002: estado = 7003;
7003: estado = 7004;
7004: estado = 7005;
7005: estado = 7006;
7006: estado = 7007;
7007: estado = 7008;
7008: estado = 7009;
7009: estado = 7010;
7010: estado = 7011;
7011: estado = 7012;
7012: estado = 7013;
7013: estado = 7014;
7014: estado = 7015;
7015: estado = 7016;
7016: estado = 7017;
7017: estado = 7018;
7018: estado = 7019;
7019: estado = 7020;
7020: estado = 7021;
7021: estado = 7022;
7022: estado = 7023;
7023: estado = 7024;
7024: estado = 7025;
7025: estado = 7026;
7026: estado = 7027;
7027: estado = 7028;
7028: estado = 7029;
7029: estado = 7030;
7030: estado = 7031;
7031: estado = 7032;
7032: estado = 7033;
7033: estado = 7034;
7034: estado = 7035;
7035: estado = 7036;
7036: estado = 7037;
7037: estado = 7038;
7038: estado = 7039;
7039: estado = 7040;
7040: estado = 7041;
7041: estado = 7042;
7042: estado = 7043;
7043: estado = 7044;
7044: estado = 7045;
7045: estado = 7046;
7046: estado = 7047;
7047: estado = 7048;
7048: estado = 7049;
7049: estado = 7050;
7050: estado = 7051;
7051: estado = 7052;
7052: estado = 7053;
7053: estado = 7054;
7054: estado = 7055;
7055: estado = 7056;
7056: estado = 7057;
7057: estado = 7058;
7058: estado = 7059;
7059: estado = 7060;
7060: estado = 7061;
7061: estado = 7062;
7062: estado = 7063;
7063: estado = 7064;
7064: estado = 7065;
7065: estado = 7066;
7066: estado = 7067;
7067: estado = 7068;
7068: estado = 7069;
7069: estado = 7070;
7070: estado = 7071;
7071: estado = 7072;
7072: estado = 7073;
7073: estado = 7074;
7074: estado = 7075;
7075: estado = 7076;
7076: estado = 7077;
7077: estado = 7078;
7078: estado = 7079;
7079: estado = 7080;
7080: estado = 7081;
7081: estado = 7082;
7082: estado = 7083;
7083: estado = 7084;
7084: estado = 7085;
7085: estado = 7086;
7086: estado = 7087;
7087: estado = 7088;
7088: estado = 7089;
7089: estado = 7090;
7090: estado = 7091;
7091: estado = 7092;
7092: estado = 7093;
7093: estado = 7094;
7094: estado = 7095;
7095: estado = 7096;
7096: estado = 7097;
7097: estado = 7098;
7098: estado = 7099;
7099: estado = 7100;
7100: estado = 7101;
7101: estado = 7102;
7102: estado = 7103;
7103: estado = 7104;
7104: estado = 7105;
7105: estado = 7106;
7106: estado = 7107;
7107: estado = 7108;
7108: estado = 7109;
7109: estado = 7110;
7110: estado = 7111;
7111: estado = 7112;
7112: estado = 7113;
7113: estado = 7114;
7114: estado = 7115;
7115: estado = 7116;
7116: estado = 7117;
7117: estado = 7118;
7118: estado = 7119;
7119: estado = 7120;
7120: estado = 7121;
7121: estado = 7122;
7122: estado = 7123;
7123: estado = 7124;
7124: estado = 7125;
7125: estado = 7126;
7126: estado = 7127;
7127: estado = 7128;
7128: estado = 7129;
7129: estado = 7130;
7130: estado = 7131;
7131: estado = 7132;
7132: estado = 7133;
7133: estado = 7134;
7134: estado = 7135;
7135: estado = 7136;
7136: estado = 7137;
7137: estado = 7138;
7138: estado = 7139;
7139: estado = 7140;
7140: estado = 7141;
7141: estado = 7142;
7142: estado = 7143;
7143: estado = 7144;
7144: estado = 7145;
7145: estado = 7146;
7146: estado = 7147;
7147: estado = 7148;
7148: estado = 7149;
7149: estado = 7150;
7150: estado = 7151;
7151: estado = 7152;
7152: estado = 7153;
7153: estado = 7154;
7154: estado = 7155;
7155: estado = 7156;
7156: estado = 7157;
7157: estado = 7158;
7158: estado = 7159;
7159: estado = 7160;
7160: estado = 7161;
7161: estado = 7162;
7162: estado = 7163;
7163: estado = 7164;
7164: estado = 7165;
7165: estado = 7166;
7166: estado = 7167;
7167: estado = 7168;
7168: estado = 7169;
7169: estado = 7170;
7170: estado = 7171;
7171: estado = 7172;
7172: estado = 7173;
7173: estado = 7174;
7174: estado = 7175;
7175: estado = 7176;
7176: estado = 7177;
7177: estado = 7178;
7178: estado = 7179;
7179: estado = 7180;
7180: estado = 7181;
7181: estado = 7182;
7182: estado = 7183;
7183: estado = 7184;
7184: estado = 7185;
7185: estado = 7186;
7186: estado = 7187;
7187: estado = 7188;
7188: estado = 7189;
7189: estado = 7190;
7190: estado = 7191;
7191: estado = 7192;
7192: estado = 7193;
7193: estado = 7194;
7194: estado = 7195;
7195: estado = 7196;
7196: estado = 7197;
7197: estado = 7198;
7198: estado = 7199;
7199: estado = 7200;
7200: estado = 7201;
7201: estado = 7202;
7202: estado = 7203;
7203: estado = 7204;
7204: estado = 7205;
7205: estado = 7206;
7206: estado = 7207;
7207: estado = 7208;
7208: estado = 7209;
7209: estado = 7210;
7210: estado = 7211;
7211: estado = 7212;
7212: estado = 7213;
7213: estado = 7214;
7214: estado = 7215;
7215: estado = 7216;
7216: estado = 7217;
7217: estado = 7218;
7218: estado = 7219;
7219: estado = 7220;
7220: estado = 7221;
7221: estado = 7222;
7222: estado = 7223;
7223: estado = 7224;
7224: estado = 7225;
7225: estado = 7226;
7226: estado = 7227;
7227: estado = 7228;
7228: estado = 7229;
7229: estado = 7230;
7230: estado = 7231;
7231: estado = 7232;
7232: estado = 7233;
7233: estado = 7234;
7234: estado = 7235;
7235: estado = 7236;
7236: estado = 7237;
7237: estado = 7238;
7238: estado = 7239;
7239: estado = 7240;
7240: estado = 7241;
7241: estado = 7242;
7242: estado = 7243;
7243: estado = 7244;
7244: estado = 7245;
7245: estado = 7246;
7246: estado = 7247;
7247: estado = 7248;
7248: estado = 7249;
7249: estado = 7250;
7250: estado = 7251;
7251: estado = 7252;
7252: estado = 7253;
7253: estado = 7254;
7254: estado = 7255;
7255: estado = 7256;
7256: estado = 7257;
7257: estado = 7258;
7258: estado = 7259;
7259: estado = 7260;
7260: estado = 7261;
7261: estado = 7262;
7262: estado = 7263;
7263: estado = 7264;
7264: estado = 7265;
7265: estado = 7266;
7266: estado = 7267;
7267: estado = 7268;
7268: estado = 7269;
7269: estado = 7270;
7270: estado = 7271;
7271: estado = 7272;
7272: estado = 7273;
7273: estado = 7274;
7274: estado = 7275;
7275: estado = 7276;
7276: estado = 7277;
7277: estado = 7278;
7278: estado = 7279;
7279: estado = 7280;
7280: estado = 7281;
7281: estado = 7282;
7282: estado = 7283;
7283: estado = 7284;
7284: estado = 7285;
7285: estado = 7286;
7286: estado = 7287;
7287: estado = 7288;
7288: estado = 7289;
7289: estado = 7290;
7290: estado = 7291;
7291: estado = 7292;
7292: estado = 7293;
7293: estado = 7294;
7294: estado = 7295;
7295: estado = 7296;
7296: estado = 7297;
7297: estado = 7298;
7298: estado = 7299;
7299: estado = 7300;
7300: estado = 7301;
7301: estado = 7302;
7302: estado = 7303;
7303: estado = 7304;
7304: estado = 7305;
7305: estado = 7306;
7306: estado = 7307;
7307: estado = 7308;
7308: estado = 7309;
7309: estado = 7310;
7310: estado = 7311;
7311: estado = 7312;
7312: estado = 7313;
7313: estado = 7314;
7314: estado = 7315;
7315: estado = 7316;
7316: estado = 7317;
7317: estado = 7318;
7318: estado = 7319;
7319: estado = 7320;
7320: estado = 7321;
7321: estado = 7322;
7322: estado = 7323;
7323: estado = 7324;
7324: estado = 7325;
7325: estado = 7326;
7326: estado = 7327;
7327: estado = 7328;
7328: estado = 7329;
7329: estado = 7330;
7330: estado = 7331;
7331: estado = 7332;
7332: estado = 7333;
7333: estado = 7334;
7334: estado = 7335;
7335: estado = 7336;
7336: estado = 7337;
7337: estado = 7338;
7338: estado = 7339;
7339: estado = 7340;
7340: estado = 7341;
7341: estado = 7342;
7342: estado = 7343;
7343: estado = 7344;
7344: estado = 7345;
7345: estado = 7346;
7346: estado = 7347;
7347: estado = 7348;
7348: estado = 7349;
7349: estado = 7350;
7350: estado = 7351;
7351: estado = 7352;
7352: estado = 7353;
7353: estado = 7354;
7354: estado = 7355;
7355: estado = 7356;
7356: estado = 7357;
7357: estado = 7358;
7358: estado = 7359;
7359: estado = 7360;
7360: estado = 7361;
7361: estado = 7362;
7362: estado = 7363;
7363: estado = 7364;
7364: estado = 7365;
7365: estado = 7366;
7366: estado = 7367;
7367: estado = 7368;
7368: estado = 7369;
7369: estado = 7370;
7370: estado = 7371;
7371: estado = 7372;
7372: estado = 7373;
7373: estado = 7374;
7374: estado = 7375;
7375: estado = 7376;
7376: estado = 7377;
7377: estado = 7378;
7378: estado = 7379;
7379: estado = 7380;
7380: estado = 7381;
7381: estado = 7382;
7382: estado = 7383;
7383: estado = 7384;
7384: estado = 7385;
7385: estado = 7386;
7386: estado = 7387;
7387: estado = 7388;
7388: estado = 7389;
7389: estado = 7390;
7390: estado = 7391;
7391: estado = 7392;
7392: estado = 7393;
7393: estado = 7394;
7394: estado = 7395;
7395: estado = 7396;
7396: estado = 7397;
7397: estado = 7398;
7398: estado = 7399;
7399: estado = 7400;
7400: estado = 7401;
7401: estado = 7402;
7402: estado = 7403;
7403: estado = 7404;
7404: estado = 7405;
7405: estado = 7406;
7406: estado = 7407;
7407: estado = 7408;
7408: estado = 7409;
7409: estado = 7410;
7410: estado = 7411;
7411: estado = 7412;
7412: estado = 7413;
7413: estado = 7414;
7414: estado = 7415;
7415: estado = 7416;
7416: estado = 7417;
7417: estado = 7418;
7418: estado = 7419;
7419: estado = 7420;
7420: estado = 7421;
7421: estado = 7422;
7422: estado = 7423;
7423: estado = 7424;
7424: estado = 7425;
7425: estado = 7426;
7426: estado = 7427;
7427: estado = 7428;
7428: estado = 7429;
7429: estado = 7430;
7430: estado = 7431;
7431: estado = 7432;
7432: estado = 7433;
7433: estado = 7434;
7434: estado = 7435;
7435: estado = 7436;
7436: estado = 7437;
7437: estado = 7438;
7438: estado = 7439;
7439: estado = 7440;
7440: estado = 7441;
7441: estado = 7442;
7442: estado = 7443;
7443: estado = 7444;
7444: estado = 7445;
7445: estado = 7446;
7446: estado = 7447;
7447: estado = 7448;
7448: estado = 7449;
7449: estado = 7450;
7450: estado = 7451;
7451: estado = 7452;
7452: estado = 7453;
7453: estado = 7454;
7454: estado = 7455;
7455: estado = 7456;
7456: estado = 7457;
7457: estado = 7458;
7458: estado = 7459;
7459: estado = 7460;
7460: estado = 7461;
7461: estado = 7462;
7462: estado = 7463;
7463: estado = 7464;
7464: estado = 7465;
7465: estado = 7466;
7466: estado = 7467;
7467: estado = 7468;
7468: estado = 7469;
7469: estado = 7470;
7470: estado = 7471;
7471: estado = 7472;
7472: estado = 7473;
7473: estado = 7474;
7474: estado = 7475;
7475: estado = 7476;
7476: estado = 7477;
7477: estado = 7478;
7478: estado = 7479;
7479: estado = 7480;
7480: estado = 7481;
7481: estado = 7482;
7482: estado = 7483;
7483: estado = 7484;
7484: estado = 7485;
7485: estado = 7486;
7486: estado = 7487;
7487: estado = 7488;
7488: estado = 7489;
7489: estado = 7490;
7490: estado = 7491;
7491: estado = 7492;
7492: estado = 7493;
7493: estado = 7494;
7494: estado = 7495;
7495: estado = 7496;
7496: estado = 7497;
7497: estado = 7498;
7498: estado = 7499;
7499: estado = 7500;
7500: estado = 7501;
7501: estado = 7502;
7502: estado = 7503;
7503: estado = 7504;
7504: estado = 7505;
7505: estado = 7506;
7506: estado = 7507;
7507: estado = 7508;
7508: estado = 7509;
7509: estado = 7510;
7510: estado = 7511;
7511: estado = 7512;
7512: estado = 7513;
7513: estado = 7514;
7514: estado = 7515;
7515: estado = 7516;
7516: estado = 7517;
7517: estado = 7518;
7518: estado = 7519;
7519: estado = 7520;
7520: estado = 7521;
7521: estado = 7522;
7522: estado = 7523;
7523: estado = 7524;
7524: estado = 7525;
7525: estado = 7526;
7526: estado = 7527;
7527: estado = 7528;
7528: estado = 7529;
7529: estado = 7530;
7530: estado = 7531;
7531: estado = 7532;
7532: estado = 7533;
7533: estado = 7534;
7534: estado = 7535;
7535: estado = 7536;
7536: estado = 7537;
7537: estado = 7538;
7538: estado = 7539;
7539: estado = 7540;
7540: estado = 7541;
7541: estado = 7542;
7542: estado = 7543;
7543: estado = 7544;
7544: estado = 7545;
7545: estado = 7546;
7546: estado = 7547;
7547: estado = 7548;
7548: estado = 7549;
7549: estado = 7550;
7550: estado = 7551;
7551: estado = 7552;
7552: estado = 7553;
7553: estado = 7554;
7554: estado = 7555;
7555: estado = 7556;
7556: estado = 7557;
7557: estado = 7558;
7558: estado = 7559;
7559: estado = 7560;
7560: estado = 7561;
7561: estado = 7562;
7562: estado = 7563;
7563: estado = 7564;
7564: estado = 7565;
7565: estado = 7566;
7566: estado = 7567;
7567: estado = 7568;
7568: estado = 7569;
7569: estado = 7570;
7570: estado = 7571;
7571: estado = 7572;
7572: estado = 7573;
7573: estado = 7574;
7574: estado = 7575;
7575: estado = 7576;
7576: estado = 7577;
7577: estado = 7578;
7578: estado = 7579;
7579: estado = 7580;
7580: estado = 7581;
7581: estado = 7582;
7582: estado = 7583;
7583: estado = 7584;
7584: estado = 7585;
7585: estado = 7586;
7586: estado = 7587;
7587: estado = 7588;
7588: estado = 7589;
7589: estado = 7590;
7590: estado = 7591;
7591: estado = 7592;
7592: estado = 7593;
7593: estado = 7594;
7594: estado = 7595;
7595: estado = 7596;
7596: estado = 7597;
7597: estado = 7598;
7598: estado = 7599;
7599: estado = 7600;
7600: estado = 7601;
7601: estado = 7602;
7602: estado = 7603;
7603: estado = 7604;
7604: estado = 7605;
7605: estado = 7606;
7606: estado = 7607;
7607: estado = 7608;
7608: estado = 7609;
7609: estado = 7610;
7610: estado = 7611;
7611: estado = 7612;
7612: estado = 7613;
7613: estado = 7614;
7614: estado = 7615;
7615: estado = 7616;
7616: estado = 7617;
7617: estado = 7618;
7618: estado = 7619;
7619: estado = 7620;
7620: estado = 7621;
7621: estado = 7622;
7622: estado = 7623;
7623: estado = 7624;
7624: estado = 7625;
7625: estado = 7626;
7626: estado = 7627;
7627: estado = 7628;
7628: estado = 7629;
7629: estado = 7630;
7630: estado = 7631;
7631: estado = 7632;
7632: estado = 7633;
7633: estado = 7634;
7634: estado = 7635;
7635: estado = 7636;
7636: estado = 7637;
7637: estado = 7638;
7638: estado = 7639;
7639: estado = 7640;
7640: estado = 7641;
7641: estado = 7642;
7642: estado = 7643;
7643: estado = 7644;
7644: estado = 7645;
7645: estado = 7646;
7646: estado = 7647;
7647: estado = 7648;
7648: estado = 7649;
7649: estado = 7650;
7650: estado = 7651;
7651: estado = 7652;
7652: estado = 7653;
7653: estado = 7654;
7654: estado = 7655;
7655: estado = 7656;
7656: estado = 7657;
7657: estado = 7658;
7658: estado = 7659;
7659: estado = 7660;
7660: estado = 7661;
7661: estado = 7662;
7662: estado = 7663;
7663: estado = 7664;
7664: estado = 7665;
7665: estado = 7666;
7666: estado = 7667;
7667: estado = 7668;
7668: estado = 7669;
7669: estado = 7670;
7670: estado = 7671;
7671: estado = 7672;
7672: estado = 7673;
7673: estado = 7674;
7674: estado = 7675;
7675: estado = 7676;
7676: estado = 7677;
7677: estado = 7678;
7678: estado = 7679;
7679: estado = 7680;
7680: estado = 7681;
7681: estado = 7682;
7682: estado = 7683;
7683: estado = 7684;
7684: estado = 7685;
7685: estado = 7686;
7686: estado = 7687;
7687: estado = 7688;
7688: estado = 7689;
7689: estado = 7690;
7690: estado = 7691;
7691: estado = 7692;
7692: estado = 7693;
7693: estado = 7694;
7694: estado = 7695;
7695: estado = 7696;
7696: estado = 7697;
7697: estado = 7698;
7698: estado = 7699;
7699: estado = 7700;
7700: estado = 7701;
7701: estado = 7702;
7702: estado = 7703;
7703: estado = 7704;
7704: estado = 7705;
7705: estado = 7706;
7706: estado = 7707;
7707: estado = 7708;
7708: estado = 7709;
7709: estado = 7710;
7710: estado = 7711;
7711: estado = 7712;
7712: estado = 7713;
7713: estado = 7714;
7714: estado = 7715;
7715: estado = 7716;
7716: estado = 7717;
7717: estado = 7718;
7718: estado = 7719;
7719: estado = 7720;
7720: estado = 7721;
7721: estado = 7722;
7722: estado = 7723;
7723: estado = 7724;
7724: estado = 7725;
7725: estado = 7726;
7726: estado = 7727;
7727: estado = 7728;
7728: estado = 7729;
7729: estado = 7730;
7730: estado = 7731;
7731: estado = 7732;
7732: estado = 7733;
7733: estado = 7734;
7734: estado = 7735;
7735: estado = 7736;
7736: estado = 7737;
7737: estado = 7738;
7738: estado = 7739;
7739: estado = 7740;
7740: estado = 7741;
7741: estado = 7742;
7742: estado = 7743;
7743: estado = 7744;
7744: estado = 7745;
7745: estado = 7746;
7746: estado = 7747;
7747: estado = 7748;
7748: estado = 7749;
7749: estado = 7750;
7750: estado = 7751;
7751: estado = 7752;
7752: estado = 7753;
7753: estado = 7754;
7754: estado = 7755;
7755: estado = 7756;
7756: estado = 7757;
7757: estado = 7758;
7758: estado = 7759;
7759: estado = 7760;
7760: estado = 7761;
7761: estado = 7762;
7762: estado = 7763;
7763: estado = 7764;
7764: estado = 7765;
7765: estado = 7766;
7766: estado = 7767;
7767: estado = 7768;
7768: estado = 7769;
7769: estado = 7770;
7770: estado = 7771;
7771: estado = 7772;
7772: estado = 7773;
7773: estado = 7774;
7774: estado = 7775;
7775: estado = 7776;
7776: estado = 7777;
7777: estado = 7778;
7778: estado = 7779;
7779: estado = 7780;
7780: estado = 7781;
7781: estado = 7782;
7782: estado = 7783;
7783: estado = 7784;
7784: estado = 7785;
7785: estado = 7786;
7786: estado = 7787;
7787: estado = 7788;
7788: estado = 7789;
7789: estado = 7790;
7790: estado = 7791;
7791: estado = 7792;
7792: estado = 7793;
7793: estado = 7794;
7794: estado = 7795;
7795: estado = 7796;
7796: estado = 7797;
7797: estado = 7798;
7798: estado = 7799;
7799: estado = 7800;
7800: estado = 7801;
7801: estado = 7802;
7802: estado = 7803;
7803: estado = 7804;
7804: estado = 7805;
7805: estado = 7806;
7806: estado = 7807;
7807: estado = 7808;
7808: estado = 7809;
7809: estado = 7810;
7810: estado = 7811;
7811: estado = 7812;
7812: estado = 7813;
7813: estado = 7814;
7814: estado = 7815;
7815: estado = 7816;
7816: estado = 7817;
7817: estado = 7818;
7818: estado = 7819;
7819: estado = 7820;
7820: estado = 7821;
7821: estado = 7822;
7822: estado = 7823;
7823: estado = 7824;
7824: estado = 7825;
7825: estado = 7826;
7826: estado = 7827;
7827: estado = 7828;
7828: estado = 7829;
7829: estado = 7830;
7830: estado = 7831;
7831: estado = 7832;
7832: estado = 7833;
7833: estado = 7834;
7834: estado = 7835;
7835: estado = 7836;
7836: estado = 7837;
7837: estado = 7838;
7838: estado = 7839;
7839: estado = 7840;
7840: estado = 7841;
7841: estado = 7842;
7842: estado = 7843;
7843: estado = 7844;
7844: estado = 7845;
7845: estado = 7846;
7846: estado = 7847;
7847: estado = 7848;
7848: estado = 7849;
7849: estado = 7850;
7850: estado = 7851;
7851: estado = 7852;
7852: estado = 7853;
7853: estado = 7854;
7854: estado = 7855;
7855: estado = 7856;
7856: estado = 7857;
7857: estado = 7858;
7858: estado = 7859;
7859: estado = 7860;
7860: estado = 7861;
7861: estado = 7862;
7862: estado = 7863;
7863: estado = 7864;
7864: estado = 7865;
7865: estado = 7866;
7866: estado = 7867;
7867: estado = 7868;
7868: estado = 7869;
7869: estado = 7870;
7870: estado = 7871;
7871: estado = 7872;
7872: estado = 7873;
7873: estado = 7874;
7874: estado = 7875;
7875: estado = 7876;
7876: estado = 7877;
7877: estado = 7878;
7878: estado = 7879;
7879: estado = 7880;
7880: estado = 7881;
7881: estado = 7882;
7882: estado = 7883;
7883: estado = 7884;
7884: estado = 7885;
7885: estado = 7886;
7886: estado = 7887;
7887: estado = 7888;
7888: estado = 7889;
7889: estado = 7890;
7890: estado = 7891;
7891: estado = 7892;
7892: estado = 7893;
7893: estado = 7894;
7894: estado = 7895;
7895: estado = 7896;
7896: estado = 7897;
7897: estado = 7898;
7898: estado = 7899;
7899: estado = 7900;
7900: estado = 7901;
7901: estado = 7902;
7902: estado = 7903;
7903: estado = 7904;
7904: estado = 7905;
7905: estado = 7906;
7906: estado = 7907;
7907: estado = 7908;
7908: estado = 7909;
7909: estado = 7910;
7910: estado = 7911;
7911: estado = 7912;
7912: estado = 7913;
7913: estado = 7914;
7914: estado = 7915;
7915: estado = 7916;
7916: estado = 7917;
7917: estado = 7918;
7918: estado = 7919;
7919: estado = 7920;
7920: estado = 7921;
7921: estado = 7922;
7922: estado = 7923;
7923: estado = 7924;
7924: estado = 7925;
7925: estado = 7926;
7926: estado = 7927;
7927: estado = 7928;
7928: estado = 7929;
7929: estado = 7930;
7930: estado = 7931;
7931: estado = 7932;
7932: estado = 7933;
7933: estado = 7934;
7934: estado = 7935;
7935: estado = 7936;
7936: estado = 7937;
7937: estado = 7938;
7938: estado = 7939;
7939: estado = 7940;
7940: estado = 7941;
7941: estado = 7942;
7942: estado = 7943;
7943: estado = 7944;
7944: estado = 7945;
7945: estado = 7946;
7946: estado = 7947;
7947: estado = 7948;
7948: estado = 7949;
7949: estado = 7950;
7950: estado = 7951;
7951: estado = 7952;
7952: estado = 7953;
7953: estado = 7954;
7954: estado = 7955;
7955: estado = 7956;
7956: estado = 7957;
7957: estado = 7958;
7958: estado = 7959;
7959: estado = 7960;
7960: estado = 7961;
7961: estado = 7962;
7962: estado = 7963;
7963: estado = 7964;
7964: estado = 7965;
7965: estado = 7966;
7966: estado = 7967;
7967: estado = 7968;
7968: estado = 7969;
7969: estado = 7970;
7970: estado = 7971;
7971: estado = 7972;
7972: estado = 7973;
7973: estado = 7974;
7974: estado = 7975;
7975: estado = 7976;
7976: estado = 7977;
7977: estado = 7978;
7978: estado = 7979;
7979: estado = 7980;
7980: estado = 7981;
7981: estado = 7982;
7982: estado = 7983;
7983: estado = 7984;
7984: estado = 7985;
7985: estado = 7986;
7986: estado = 7987;
7987: estado = 7988;
7988: estado = 7989;
7989: estado = 7990;
7990: estado = 7991;
7991: estado = 7992;
7992: estado = 7993;
7993: estado = 7994;
7994: estado = 7995;
7995: estado = 7996;
7996: estado = 7997;
7997: estado = 7998;
7998: estado = 7999;
7999: estado = 8000;
8000: estado = 8001;
8001: estado = 8002;
8002: estado = 8003;
8003: estado = 8004;
8004: estado = 8005;
8005: estado = 8006;
8006: estado = 8007;
8007: estado = 8008;
8008: estado = 8009;
8009: estado = 8010;
8010: estado = 8011;
8011: estado = 8012;
8012: estado = 8013;
8013: estado = 8014;
8014: estado = 8015;
8015: estado = 8016;
8016: estado = 8017;
8017: estado = 8018;
8018: estado = 8019;
8019: estado = 8020;
8020: estado = 8021;
8021: estado = 8022;
8022: estado = 8023;
8023: estado = 8024;
8024: estado = 8025;
8025: estado = 8026;
8026: estado = 8027;
8027: estado = 8028;
8028: estado = 8029;
8029: estado = 8030;
8030: estado = 8031;
8031: estado = 8032;
8032: estado = 8033;
8033: estado = 8034;
8034: estado = 8035;
8035: estado = 8036;
8036: estado = 8037;
8037: estado = 8038;
8038: estado = 8039;
8039: estado = 8040;
8040: estado = 8041;
8041: estado = 8042;
8042: estado = 8043;
8043: estado = 8044;
8044: estado = 8045;
8045: estado = 8046;
8046: estado = 8047;
8047: estado = 8048;
8048: estado = 8049;
8049: estado = 8050;
8050: estado = 8051;
8051: estado = 8052;
8052: estado = 8053;
8053: estado = 8054;
8054: estado = 8055;
8055: estado = 8056;
8056: estado = 8057;
8057: estado = 8058;
8058: estado = 8059;
8059: estado = 8060;
8060: estado = 8061;
8061: estado = 8062;
8062: estado = 8063;
8063: estado = 8064;
8064: estado = 8065;
8065: estado = 8066;
8066: estado = 8067;
8067: estado = 8068;
8068: estado = 8069;
8069: estado = 8070;
8070: estado = 8071;
8071: estado = 8072;
8072: estado = 8073;
8073: estado = 8074;
8074: estado = 8075;
8075: estado = 8076;
8076: estado = 8077;
8077: estado = 8078;
8078: estado = 8079;
8079: estado = 8080;
8080: estado = 8081;
8081: estado = 8082;
8082: estado = 8083;
8083: estado = 8084;
8084: estado = 8085;
8085: estado = 8086;
8086: estado = 8087;
8087: estado = 8088;
8088: estado = 8089;
8089: estado = 8090;
8090: estado = 8091;
8091: estado = 8092;
8092: estado = 8093;
8093: estado = 8094;
8094: estado = 8095;
8095: estado = 8096;
8096: estado = 8097;
8097: estado = 8098;
8098: estado = 8099;
8099: estado = 8100;
8100: estado = 8101;
8101: estado = 8102;
8102: estado = 8103;
8103: estado = 8104;
8104: estado = 8105;
8105: estado = 8106;
8106: estado = 8107;
8107: estado = 8108;
8108: estado = 8109;
8109: estado = 8110;
8110: estado = 8111;
8111: estado = 8112;
8112: estado = 8113;
8113: estado = 8114;
8114: estado = 8115;
8115: estado = 8116;
8116: estado = 8117;
8117: estado = 8118;
8118: estado = 8119;
8119: estado = 8120;
8120: estado = 8121;
8121: estado = 8122;
8122: estado = 8123;
8123: estado = 8124;
8124: estado = 8125;
8125: estado = 8126;
8126: estado = 8127;
8127: estado = 8128;
8128: estado = 8129;
8129: estado = 8130;
8130: estado = 8131;
8131: estado = 8132;
8132: estado = 8133;
8133: estado = 8134;
8134: estado = 8135;
8135: estado = 8136;
8136: estado = 8137;
8137: estado = 8138;
8138: estado = 8139;
8139: estado = 8140;
8140: estado = 8141;
8141: estado = 8142;
8142: estado = 8143;
8143: estado = 8144;
8144: estado = 8145;
8145: estado = 8146;
8146: estado = 8147;
8147: estado = 8148;
8148: estado = 8149;
8149: estado = 8150;
8150: estado = 8151;
8151: estado = 8152;
8152: estado = 8153;
8153: estado = 8154;
8154: estado = 8155;
8155: estado = 8156;
8156: estado = 8157;
8157: estado = 8158;
8158: estado = 8159;
8159: estado = 8160;
8160: estado = 8161;
8161: estado = 8162;
8162: estado = 8163;
8163: estado = 8164;
8164: estado = 8165;
8165: estado = 8166;
8166: estado = 8167;
8167: estado = 8168;
8168: estado = 8169;
8169: estado = 8170;
8170: estado = 8171;
8171: estado = 8172;
8172: estado = 8173;
8173: estado = 8174;
8174: estado = 8175;
8175: estado = 8176;
8176: estado = 8177;
8177: estado = 8178;
8178: estado = 8179;
8179: estado = 8180;
8180: estado = 8181;
8181: estado = 8182;
8182: estado = 8183;
8183: estado = 8184;
8184: estado = 8185;
8185: estado = 8186;
8186: estado = 8187;
8187: estado = 8188;
8188: estado = 8189;
8189: estado = 8190;
8190: estado = 8191;
8191: estado = 8192;
8192: estado = 8193;
8193: estado = 8194;
8194: estado = 8195;
8195: estado = 8196;
8196: estado = 8197;
8197: estado = 8198;
8198: estado = 8199;
8199: estado = 8200;
8200: estado = 8201;
8201: estado = 8202;
8202: estado = 8203;
8203: estado = 8204;
8204: estado = 8205;
8205: estado = 8206;
8206: estado = 8207;
8207: estado = 8208;
8208: estado = 8209;
8209: estado = 8210;
8210: estado = 8211;
8211: estado = 8212;
8212: estado = 8213;
8213: estado = 8214;
8214: estado = 8215;
8215: estado = 8216;
8216: estado = 8217;
8217: estado = 8218;
8218: estado = 8219;
8219: estado = 8220;
8220: estado = 8221;
8221: estado = 8222;
8222: estado = 8223;
8223: estado = 8224;
8224: estado = 8225;
8225: estado = 8226;
8226: estado = 8227;
8227: estado = 8228;
8228: estado = 8229;
8229: estado = 8230;
8230: estado = 8231;
8231: estado = 8232;
8232: estado = 8233;
8233: estado = 8234;
8234: estado = 8235;
8235: estado = 8236;
8236: estado = 8237;
8237: estado = 8238;
8238: estado = 8239;
8239: estado = 8240;
8240: estado = 8241;
8241: estado = 8242;
8242: estado = 8243;
8243: estado = 8244;
8244: estado = 8245;
8245: estado = 8246;
8246: estado = 8247;
8247: estado = 8248;
8248: estado = 8249;
8249: estado = 8250;
8250: estado = 8251;
8251: estado = 8252;
8252: estado = 8253;
8253: estado = 8254;
8254: estado = 8255;
8255: estado = 8256;
8256: estado = 8257;
8257: estado = 8258;
8258: estado = 8259;
8259: estado = 8260;
8260: estado = 8261;
8261: estado = 8262;
8262: estado = 8263;
8263: estado = 8264;
8264: estado = 8265;
8265: estado = 8266;
8266: estado = 8267;
8267: estado = 8268;
8268: estado = 8269;
8269: estado = 8270;
8270: estado = 8271;
8271: estado = 8272;
8272: estado = 8273;
8273: estado = 8274;
8274: estado = 8275;
8275: estado = 8276;
8276: estado = 8277;
8277: estado = 8278;
8278: estado = 8279;
8279: estado = 8280;
8280: estado = 8281;
8281: estado = 8282;
8282: estado = 8283;
8283: estado = 8284;
8284: estado = 8285;
8285: estado = 8286;
8286: estado = 8287;
8287: estado = 8288;
8288: estado = 8289;
8289: estado = 8290;
8290: estado = 8291;
8291: estado = 8292;
8292: estado = 8293;
8293: estado = 8294;
8294: estado = 8295;
8295: estado = 8296;
8296: estado = 8297;
8297: estado = 8298;
8298: estado = 8299;
8299: estado = 8300;
8300: estado = 8301;
8301: estado = 8302;
8302: estado = 8303;
8303: estado = 8304;
8304: estado = 8305;
8305: estado = 8306;
8306: estado = 8307;
8307: estado = 8308;
8308: estado = 8309;
8309: estado = 8310;
8310: estado = 8311;
8311: estado = 8312;
8312: estado = 8313;
8313: estado = 8314;
8314: estado = 8315;
8315: estado = 8316;
8316: estado = 8317;
8317: estado = 8318;
8318: estado = 8319;
8319: estado = 8320;
8320: estado = 8321;
8321: estado = 8322;
8322: estado = 8323;
8323: estado = 8324;
8324: estado = 8325;
8325: estado = 8326;
8326: estado = 8327;
8327: estado = 8328;
8328: estado = 8329;
8329: estado = 8330;
8330: estado = 8331;
8331: estado = 8332;
8332: estado = 8333;
8333: estado = 8334;
8334: estado = 8335;
8335: estado = 8336;
8336: estado = 8337;
8337: estado = 8338;
8338: estado = 8339;
8339: estado = 8340;
8340: estado = 8341;
8341: estado = 8342;
8342: estado = 8343;
8343: estado = 8344;
8344: estado = 8345;
8345: estado = 8346;
8346: estado = 8347;
8347: estado = 8348;
8348: estado = 8349;
8349: estado = 8350;
8350: estado = 8351;
8351: estado = 8352;
8352: estado = 8353;
8353: estado = 8354;
8354: estado = 8355;
8355: estado = 8356;
8356: estado = 8357;
8357: estado = 8358;
8358: estado = 8359;
8359: estado = 8360;
8360: estado = 8361;
8361: estado = 8362;
8362: estado = 8363;
8363: estado = 8364;
8364: estado = 8365;
8365: estado = 8366;
8366: estado = 8367;
8367: estado = 8368;
8368: estado = 8369;
8369: estado = 8370;
8370: estado = 8371;
8371: estado = 8372;
8372: estado = 8373;
8373: estado = 8374;
8374: estado = 8375;
8375: estado = 8376;
8376: estado = 8377;
8377: estado = 8378;
8378: estado = 8379;
8379: estado = 8380;
8380: estado = 8381;
8381: estado = 8382;
8382: estado = 8383;
8383: estado = 8384;
8384: estado = 8385;
8385: estado = 8386;
8386: estado = 8387;
8387: estado = 8388;
8388: estado = 8389;
8389: estado = 8390;
8390: estado = 8391;
8391: estado = 8392;
8392: estado = 8393;
8393: estado = 8394;
8394: estado = 8395;
8395: estado = 8396;
8396: estado = 8397;
8397: estado = 8398;
8398: estado = 8399;
8399: estado = 8400;
8400: estado = 8401;
8401: estado = 8402;
8402: estado = 8403;
8403: estado = 8404;
8404: estado = 8405;
8405: estado = 8406;
8406: estado = 8407;
8407: estado = 8408;
8408: estado = 8409;
8409: estado = 8410;
8410: estado = 8411;
8411: estado = 8412;
8412: estado = 8413;
8413: estado = 8414;
8414: estado = 8415;
8415: estado = 8416;
8416: estado = 8417;
8417: estado = 8418;
8418: estado = 8419;
8419: estado = 8420;
8420: estado = 8421;
8421: estado = 8422;
8422: estado = 8423;
8423: estado = 8424;
8424: estado = 8425;
8425: estado = 8426;
8426: estado = 8427;
8427: estado = 8428;
8428: estado = 8429;
8429: estado = 8430;
8430: estado = 8431;
8431: estado = 8432;
8432: estado = 8433;
8433: estado = 8434;
8434: estado = 8435;
8435: estado = 8436;
8436: estado = 8437;
8437: estado = 8438;
8438: estado = 8439;
8439: estado = 8440;
8440: estado = 8441;
8441: estado = 8442;
8442: estado = 8443;
8443: estado = 8444;
8444: estado = 8445;
8445: estado = 8446;
8446: estado = 8447;
8447: estado = 8448;
8448: estado = 8449;
8449: estado = 8450;
8450: estado = 8451;
8451: estado = 8452;
8452: estado = 8453;
8453: estado = 8454;
8454: estado = 8455;
8455: estado = 8456;
8456: estado = 8457;
8457: estado = 8458;
8458: estado = 8459;
8459: estado = 8460;
8460: estado = 8461;
8461: estado = 8462;
8462: estado = 8463;
8463: estado = 8464;
8464: estado = 8465;
8465: estado = 8466;
8466: estado = 8467;
8467: estado = 8468;
8468: estado = 8469;
8469: estado = 8470;
8470: estado = 8471;
8471: estado = 8472;
8472: estado = 8473;
8473: estado = 8474;
8474: estado = 8475;
8475: estado = 8476;
8476: estado = 8477;
8477: estado = 8478;
8478: estado = 8479;
8479: estado = 8480;
8480: estado = 8481;
8481: estado = 8482;
8482: estado = 8483;
8483: estado = 8484;
8484: estado = 8485;
8485: estado = 8486;
8486: estado = 8487;
8487: estado = 8488;
8488: estado = 8489;
8489: estado = 8490;
8490: estado = 8491;
8491: estado = 8492;
8492: estado = 8493;
8493: estado = 8494;
8494: estado = 8495;
8495: estado = 8496;
8496: estado = 8497;
8497: estado = 8498;
8498: estado = 8499;
8499: estado = 8500;
8500: estado = 8501;
8501: estado = 8502;
8502: estado = 8503;
8503: estado = 8504;
8504: estado = 8505;
8505: estado = 8506;
8506: estado = 8507;
8507: estado = 8508;
8508: estado = 8509;
8509: estado = 8510;
8510: estado = 8511;
8511: estado = 8512;
8512: estado = 8513;
8513: estado = 8514;
8514: estado = 8515;
8515: estado = 8516;
8516: estado = 8517;
8517: estado = 8518;
8518: estado = 8519;
8519: estado = 8520;
8520: estado = 8521;
8521: estado = 8522;
8522: estado = 8523;
8523: estado = 8524;
8524: estado = 8525;
8525: estado = 8526;
8526: estado = 8527;
8527: estado = 8528;
8528: estado = 8529;
8529: estado = 8530;
8530: estado = 8531;
8531: estado = 8532;
8532: estado = 8533;
8533: estado = 8534;
8534: estado = 8535;
8535: estado = 8536;
8536: estado = 8537;
8537: estado = 8538;
8538: estado = 8539;
8539: estado = 8540;
8540: estado = 8541;
8541: estado = 8542;
8542: estado = 8543;
8543: estado = 8544;
8544: estado = 8545;
8545: estado = 8546;
8546: estado = 8547;
8547: estado = 8548;
8548: estado = 8549;
8549: estado = 8550;
8550: estado = 8551;
8551: estado = 8552;
8552: estado = 8553;
8553: estado = 8554;
8554: estado = 8555;
8555: estado = 8556;
8556: estado = 8557;
8557: estado = 8558;
8558: estado = 8559;
8559: estado = 8560;
8560: estado = 8561;
8561: estado = 8562;
8562: estado = 8563;
8563: estado = 8564;
8564: estado = 8565;
8565: estado = 8566;
8566: estado = 8567;
8567: estado = 8568;
8568: estado = 8569;
8569: estado = 8570;
8570: estado = 8571;
8571: estado = 8572;
8572: estado = 8573;
8573: estado = 8574;
8574: estado = 8575;
8575: estado = 8576;
8576: estado = 8577;
8577: estado = 8578;
8578: estado = 8579;
8579: estado = 8580;
8580: estado = 8581;
8581: estado = 8582;
8582: estado = 8583;
8583: estado = 8584;
8584: estado = 8585;
8585: estado = 8586;
8586: estado = 8587;
8587: estado = 8588;
8588: estado = 8589;
8589: estado = 8590;
8590: estado = 8591;
8591: estado = 8592;
8592: estado = 8593;
8593: estado = 8594;
8594: estado = 8595;
8595: estado = 8596;
8596: estado = 8597;
8597: estado = 8598;
8598: estado = 8599;
8599: estado = 8600;
8600: estado = 8601;
8601: estado = 8602;
8602: estado = 8603;
8603: estado = 8604;
8604: estado = 8605;
8605: estado = 8606;
8606: estado = 8607;
8607: estado = 8608;
8608: estado = 8609;
8609: estado = 8610;
8610: estado = 8611;
8611: estado = 8612;
8612: estado = 8613;
8613: estado = 8614;
8614: estado = 8615;
8615: estado = 8616;
8616: estado = 8617;
8617: estado = 8618;
8618: estado = 8619;
8619: estado = 8620;
8620: estado = 8621;
8621: estado = 8622;
8622: estado = 8623;
8623: estado = 8624;
8624: estado = 8625;
8625: estado = 8626;
8626: estado = 8627;
8627: estado = 8628;
8628: estado = 8629;
8629: estado = 8630;
8630: estado = 8631;
8631: estado = 8632;
8632: estado = 8633;
8633: estado = 8634;
8634: estado = 8635;
8635: estado = 8636;
8636: estado = 8637;
8637: estado = 8638;
8638: estado = 8639;
8639: estado = 8640;
8640: estado = 8641;
8641: estado = 8642;
8642: estado = 8643;
8643: estado = 8644;
8644: estado = 8645;
8645: estado = 8646;
8646: estado = 8647;
8647: estado = 8648;
8648: estado = 8649;
8649: estado = 8650;
8650: estado = 8651;
8651: estado = 8652;
8652: estado = 8653;
8653: estado = 8654;
8654: estado = 8655;
8655: estado = 8656;
8656: estado = 8657;
8657: estado = 8658;
8658: estado = 8659;
8659: estado = 8660;
8660: estado = 8661;
8661: estado = 8662;
8662: estado = 8663;
8663: estado = 8664;
8664: estado = 8665;
8665: estado = 8666;
8666: estado = 8667;
8667: estado = 8668;
8668: estado = 8669;
8669: estado = 8670;
8670: estado = 8671;
8671: estado = 8672;
8672: estado = 8673;
8673: estado = 8674;
8674: estado = 8675;
8675: estado = 8676;
8676: estado = 8677;
8677: estado = 8678;
8678: estado = 8679;
8679: estado = 8680;
8680: estado = 8681;
8681: estado = 8682;
8682: estado = 8683;
8683: estado = 8684;
8684: estado = 8685;
8685: estado = 8686;
8686: estado = 8687;
8687: estado = 8688;
8688: estado = 8689;
8689: estado = 8690;
8690: estado = 8691;
8691: estado = 8692;
8692: estado = 8693;
8693: estado = 8694;
8694: estado = 8695;
8695: estado = 8696;
8696: estado = 8697;
8697: estado = 8698;
8698: estado = 8699;
8699: estado = 8700;
8700: estado = 8701;
8701: estado = 8702;
8702: estado = 8703;
8703: estado = 8704;
8704: estado = 8705;
8705: estado = 8706;
8706: estado = 8707;
8707: estado = 8708;
8708: estado = 8709;
8709: estado = 8710;
8710: estado = 8711;
8711: estado = 8712;
8712: estado = 8713;
8713: estado = 8714;
8714: estado = 8715;
8715: estado = 8716;
8716: estado = 8717;
8717: estado = 8718;
8718: estado = 8719;
8719: estado = 8720;
8720: estado = 8721;
8721: estado = 8722;
8722: estado = 8723;
8723: estado = 8724;
8724: estado = 8725;
8725: estado = 8726;
8726: estado = 8727;
8727: estado = 8728;
8728: estado = 8729;
8729: estado = 8730;
8730: estado = 8731;
8731: estado = 8732;
8732: estado = 8733;
8733: estado = 8734;
8734: estado = 8735;
8735: estado = 8736;
8736: estado = 8737;
8737: estado = 8738;
8738: estado = 8739;
8739: estado = 8740;
8740: estado = 8741;
8741: estado = 8742;
8742: estado = 8743;
8743: estado = 8744;
8744: estado = 8745;
8745: estado = 8746;
8746: estado = 8747;
8747: estado = 8748;
8748: estado = 8749;
8749: estado = 8750;
8750: estado = 8751;
8751: estado = 8752;
8752: estado = 8753;
8753: estado = 8754;
8754: estado = 8755;
8755: estado = 8756;
8756: estado = 8757;
8757: estado = 8758;
8758: estado = 8759;
8759: estado = 8760;
8760: estado = 8761;
8761: estado = 8762;
8762: estado = 8763;
8763: estado = 8764;
8764: estado = 8765;
8765: estado = 8766;
8766: estado = 8767;
8767: estado = 8768;
8768: estado = 8769;
8769: estado = 8770;
8770: estado = 8771;
8771: estado = 8772;
8772: estado = 8773;
8773: estado = 8774;
8774: estado = 8775;
8775: estado = 8776;
8776: estado = 8777;
8777: estado = 8778;
8778: estado = 8779;
8779: estado = 8780;
8780: estado = 8781;
8781: estado = 8782;
8782: estado = 8783;
8783: estado = 8784;
8784: estado = 8785;
8785: estado = 8786;
8786: estado = 8787;
8787: estado = 8788;
8788: estado = 8789;
8789: estado = 8790;
8790: estado = 8791;
8791: estado = 8792;
8792: estado = 8793;
8793: estado = 8794;
8794: estado = 8795;
8795: estado = 8796;
8796: estado = 8797;
8797: estado = 8798;
8798: estado = 8799;
8799: estado = 8800;
8800: estado = 8801;
8801: estado = 8802;
8802: estado = 8803;
8803: estado = 8804;
8804: estado = 8805;
8805: estado = 8806;
8806: estado = 8807;
8807: estado = 8808;
8808: estado = 8809;
8809: estado = 8810;
8810: estado = 8811;
8811: estado = 8812;
8812: estado = 8813;
8813: estado = 8814;
8814: estado = 8815;
8815: estado = 8816;
8816: estado = 8817;
8817: estado = 8818;
8818: estado = 8819;
8819: estado = 8820;
8820: estado = 8821;
8821: estado = 8822;
8822: estado = 8823;
8823: estado = 8824;
8824: estado = 8825;
8825: estado = 8826;
8826: estado = 8827;
8827: estado = 8828;
8828: estado = 8829;
8829: estado = 8830;
8830: estado = 8831;
8831: estado = 8832;
8832: estado = 8833;
8833: estado = 8834;
8834: estado = 8835;
8835: estado = 8836;
8836: estado = 8837;
8837: estado = 8838;
8838: estado = 8839;
8839: estado = 8840;
8840: estado = 8841;
8841: estado = 8842;
8842: estado = 8843;
8843: estado = 8844;
8844: estado = 8845;
8845: estado = 8846;
8846: estado = 8847;
8847: estado = 8848;
8848: estado = 8849;
8849: estado = 8850;
8850: estado = 8851;
8851: estado = 8852;
8852: estado = 8853;
8853: estado = 8854;
8854: estado = 8855;
8855: estado = 8856;
8856: estado = 8857;
8857: estado = 8858;
8858: estado = 8859;
8859: estado = 8860;
8860: estado = 8861;
8861: estado = 8862;
8862: estado = 8863;
8863: estado = 8864;
8864: estado = 8865;
8865: estado = 8866;
8866: estado = 8867;
8867: estado = 8868;
8868: estado = 8869;
8869: estado = 8870;
8870: estado = 8871;
8871: estado = 8872;
8872: estado = 8873;
8873: estado = 8874;
8874: estado = 8875;
8875: estado = 8876;
8876: estado = 8877;
8877: estado = 8878;
8878: estado = 8879;
8879: estado = 8880;
8880: estado = 8881;
8881: estado = 8882;
8882: estado = 8883;
8883: estado = 8884;
8884: estado = 8885;
8885: estado = 8886;
8886: estado = 8887;
8887: estado = 8888;
8888: estado = 8889;
8889: estado = 8890;
8890: estado = 8891;
8891: estado = 8892;
8892: estado = 8893;
8893: estado = 8894;
8894: estado = 8895;
8895: estado = 8896;
8896: estado = 8897;
8897: estado = 8898;
8898: estado = 8899;
8899: estado = 8900;
8900: estado = 8901;
8901: estado = 8902;
8902: estado = 8903;
8903: estado = 8904;
8904: estado = 8905;
8905: estado = 8906;
8906: estado = 8907;
8907: estado = 8908;
8908: estado = 8909;
8909: estado = 8910;
8910: estado = 8911;
8911: estado = 8912;
8912: estado = 8913;
8913: estado = 8914;
8914: estado = 8915;
8915: estado = 8916;
8916: estado = 8917;
8917: estado = 8918;
8918: estado = 8919;
8919: estado = 8920;
8920: estado = 8921;
8921: estado = 8922;
8922: estado = 8923;
8923: estado = 8924;
8924: estado = 8925;
8925: estado = 8926;
8926: estado = 8927;
8927: estado = 8928;
8928: estado = 8929;
8929: estado = 8930;
8930: estado = 8931;
8931: estado = 8932;
8932: estado = 8933;
8933: estado = 8934;
8934: estado = 8935;
8935: estado = 8936;
8936: estado = 8937;
8937: estado = 8938;
8938: estado = 8939;
8939: estado = 8940;
8940: estado = 8941;
8941: estado = 8942;
8942: estado = 8943;
8943: estado = 8944;
8944: estado = 8945;
8945: estado = 8946;
8946: estado = 8947;
8947: estado = 8948;
8948: estado = 8949;
8949: estado = 8950;
8950: estado = 8951;
8951: estado = 8952;
8952: estado = 8953;
8953: estado = 8954;
8954: estado = 8955;
8955: estado = 8956;
8956: estado = 8957;
8957: estado = 8958;
8958: estado = 8959;
8959: estado = 8960;
8960: estado = 8961;
8961: estado = 8962;
8962: estado = 8963;
8963: estado = 8964;
8964: estado = 8965;
8965: estado = 8966;
8966: estado = 8967;
8967: estado = 8968;
8968: estado = 8969;
8969: estado = 8970;
8970: estado = 8971;
8971: estado = 8972;
8972: estado = 8973;
8973: estado = 8974;
8974: estado = 8975;
8975: estado = 8976;
8976: estado = 8977;
8977: estado = 8978;
8978: estado = 8979;
8979: estado = 8980;
8980: estado = 8981;
8981: estado = 8982;
8982: estado = 8983;
8983: estado = 8984;
8984: estado = 8985;
8985: estado = 8986;
8986: estado = 8987;
8987: estado = 8988;
8988: estado = 8989;
8989: estado = 8990;
8990: estado = 8991;
8991: estado = 8992;
8992: estado = 8993;
8993: estado = 8994;
8994: estado = 8995;
8995: estado = 8996;
8996: estado = 8997;
8997: estado = 8998;
8998: estado = 8999;
8999: estado = 9000;
9000: estado = 9001;
9001: estado = 9002;
9002: estado = 9003;
9003: estado = 9004;
9004: estado = 9005;
9005: estado = 9006;
9006: estado = 9007;
9007: estado = 9008;
9008: estado = 9009;
9009: estado = 9010;
9010: estado = 9011;
9011: estado = 9012;
9012: estado = 9013;
9013: estado = 9014;
9014: estado = 9015;
9015: estado = 9016;
9016: estado = 9017;
9017: estado = 9018;
9018: estado = 9019;
9019: estado = 9020;
9020: estado = 9021;
9021: estado = 9022;
9022: estado = 9023;
9023: estado = 9024;
9024: estado = 9025;
9025: estado = 9026;
9026: estado = 9027;
9027: estado = 9028;
9028: estado = 9029;
9029: estado = 9030;
9030: estado = 9031;
9031: estado = 9032;
9032: estado = 9033;
9033: estado = 9034;
9034: estado = 9035;
9035: estado = 9036;
9036: estado = 9037;
9037: estado = 9038;
9038: estado = 9039;
9039: estado = 9040;
9040: estado = 9041;
9041: estado = 9042;
9042: estado = 9043;
9043: estado = 9044;
9044: estado = 9045;
9045: estado = 9046;
9046: estado = 9047;
9047: estado = 9048;
9048: estado = 9049;
9049: estado = 9050;
9050: estado = 9051;
9051: estado = 9052;
9052: estado = 9053;
9053: estado = 9054;
9054: estado = 9055;
9055: estado = 9056;
9056: estado = 9057;
9057: estado = 9058;
9058: estado = 9059;
9059: estado = 9060;
9060: estado = 9061;
9061: estado = 9062;
9062: estado = 9063;
9063: estado = 9064;
9064: estado = 9065;
9065: estado = 9066;
9066: estado = 9067;
9067: estado = 9068;
9068: estado = 9069;
9069: estado = 9070;
9070: estado = 9071;
9071: estado = 9072;
9072: estado = 9073;
9073: estado = 9074;
9074: estado = 9075;
9075: estado = 9076;
9076: estado = 9077;
9077: estado = 9078;
9078: estado = 9079;
9079: estado = 9080;
9080: estado = 9081;
9081: estado = 9082;
9082: estado = 9083;
9083: estado = 9084;
9084: estado = 9085;
9085: estado = 9086;
9086: estado = 9087;
9087: estado = 9088;
9088: estado = 9089;
9089: estado = 9090;
9090: estado = 9091;
9091: estado = 9092;
9092: estado = 9093;
9093: estado = 9094;
9094: estado = 9095;
9095: estado = 9096;
9096: estado = 9097;
9097: estado = 9098;
9098: estado = 9099;
9099: estado = 9100;
9100: estado = 9101;
9101: estado = 9102;
9102: estado = 9103;
9103: estado = 9104;
9104: estado = 9105;
9105: estado = 9106;
9106: estado = 9107;
9107: estado = 9108;
9108: estado = 9109;
9109: estado = 9110;
9110: estado = 9111;
9111: estado = 9112;
9112: estado = 9113;
9113: estado = 9114;
9114: estado = 9115;
9115: estado = 9116;
9116: estado = 9117;
9117: estado = 9118;
9118: estado = 9119;
9119: estado = 9120;
9120: estado = 9121;
9121: estado = 9122;
9122: estado = 9123;
9123: estado = 9124;
9124: estado = 9125;
9125: estado = 9126;
9126: estado = 9127;
9127: estado = 9128;
9128: estado = 9129;
9129: estado = 9130;
9130: estado = 9131;
9131: estado = 9132;
9132: estado = 9133;
9133: estado = 9134;
9134: estado = 9135;
9135: estado = 9136;
9136: estado = 9137;
9137: estado = 9138;
9138: estado = 9139;
9139: estado = 9140;
9140: estado = 9141;
9141: estado = 9142;
9142: estado = 9143;
9143: estado = 9144;
9144: estado = 9145;
9145: estado = 9146;
9146: estado = 9147;
9147: estado = 9148;
9148: estado = 9149;
9149: estado = 9150;
9150: estado = 9151;
9151: estado = 9152;
9152: estado = 9153;
9153: estado = 9154;
9154: estado = 9155;
9155: estado = 9156;
9156: estado = 9157;
9157: estado = 9158;
9158: estado = 9159;
9159: estado = 9160;
9160: estado = 9161;
9161: estado = 9162;
9162: estado = 9163;
9163: estado = 9164;
9164: estado = 9165;
9165: estado = 9166;
9166: estado = 9167;
9167: estado = 9168;
9168: estado = 9169;
9169: estado = 9170;
9170: estado = 9171;
9171: estado = 9172;
9172: estado = 9173;
9173: estado = 9174;
9174: estado = 9175;
9175: estado = 9176;
9176: estado = 9177;
9177: estado = 9178;
9178: estado = 9179;
9179: estado = 9180;
9180: estado = 9181;
9181: estado = 9182;
9182: estado = 9183;
9183: estado = 9184;
9184: estado = 9185;
9185: estado = 9186;
9186: estado = 9187;
9187: estado = 9188;
9188: estado = 9189;
9189: estado = 9190;
9190: estado = 9191;
9191: estado = 9192;
9192: estado = 9193;
9193: estado = 9194;
9194: estado = 9195;
9195: estado = 9196;
9196: estado = 9197;
9197: estado = 9198;
9198: estado = 9199;
9199: estado = 9200;
9200: estado = 9201;
9201: estado = 9202;
9202: estado = 9203;
9203: estado = 9204;
9204: estado = 9205;
9205: estado = 9206;
9206: estado = 9207;
9207: estado = 9208;
9208: estado = 9209;
9209: estado = 9210;
9210: estado = 9211;
9211: estado = 9212;
9212: estado = 9213;
9213: estado = 9214;
9214: estado = 9215;
9215: estado = 9216;
9216: estado = 9217;
9217: estado = 9218;
9218: estado = 9219;
9219: estado = 9220;
9220: estado = 9221;
9221: estado = 9222;
9222: estado = 9223;
9223: estado = 9224;
9224: estado = 9225;
9225: estado = 9226;
9226: estado = 9227;
9227: estado = 9228;
9228: estado = 9229;
9229: estado = 9230;
9230: estado = 9231;
9231: estado = 9232;
9232: estado = 9233;
9233: estado = 9234;
9234: estado = 9235;
9235: estado = 9236;
9236: estado = 9237;
9237: estado = 9238;
9238: estado = 9239;
9239: estado = 9240;
9240: estado = 9241;
9241: estado = 9242;
9242: estado = 9243;
9243: estado = 9244;
9244: estado = 9245;
9245: estado = 9246;
9246: estado = 9247;
9247: estado = 9248;
9248: estado = 9249;
9249: estado = 9250;
9250: estado = 9251;
9251: estado = 9252;
9252: estado = 9253;
9253: estado = 9254;
9254: estado = 9255;
9255: estado = 9256;
9256: estado = 9257;
9257: estado = 9258;
9258: estado = 9259;
9259: estado = 9260;
9260: estado = 9261;
9261: estado = 9262;
9262: estado = 9263;
9263: estado = 9264;
9264: estado = 9265;
9265: estado = 9266;
9266: estado = 9267;
9267: estado = 9268;
9268: estado = 9269;
9269: estado = 9270;
9270: estado = 9271;
9271: estado = 9272;
9272: estado = 9273;
9273: estado = 9274;
9274: estado = 9275;
9275: estado = 9276;
9276: estado = 9277;
9277: estado = 9278;
9278: estado = 9279;
9279: estado = 9280;
9280: estado = 9281;
9281: estado = 9282;
9282: estado = 9283;
9283: estado = 9284;
9284: estado = 9285;
9285: estado = 9286;
9286: estado = 9287;
9287: estado = 9288;
9288: estado = 9289;
9289: estado = 9290;
9290: estado = 9291;
9291: estado = 9292;
9292: estado = 9293;
9293: estado = 9294;
9294: estado = 9295;
9295: estado = 9296;
9296: estado = 9297;
9297: estado = 9298;
9298: estado = 9299;
9299: estado = 9300;
9300: estado = 9301;
9301: estado = 9302;
9302: estado = 9303;
9303: estado = 9304;
9304: estado = 9305;
9305: estado = 9306;
9306: estado = 9307;
9307: estado = 9308;
9308: estado = 9309;
9309: estado = 9310;
9310: estado = 9311;
9311: estado = 9312;
9312: estado = 9313;
9313: estado = 9314;
9314: estado = 9315;
9315: estado = 9316;
9316: estado = 9317;
9317: estado = 9318;
9318: estado = 9319;
9319: estado = 9320;
9320: estado = 9321;
9321: estado = 9322;
9322: estado = 9323;
9323: estado = 9324;
9324: estado = 9325;
9325: estado = 9326;
9326: estado = 9327;
9327: estado = 9328;
9328: estado = 9329;
9329: estado = 9330;
9330: estado = 9331;
9331: estado = 9332;
9332: estado = 9333;
9333: estado = 9334;
9334: estado = 9335;
9335: estado = 9336;
9336: estado = 9337;
9337: estado = 9338;
9338: estado = 9339;
9339: estado = 9340;
9340: estado = 9341;
9341: estado = 9342;
9342: estado = 9343;
9343: estado = 9344;
9344: estado = 9345;
9345: estado = 9346;
9346: estado = 9347;
9347: estado = 9348;
9348: estado = 9349;
9349: estado = 9350;
9350: estado = 9351;
9351: estado = 9352;
9352: estado = 9353;
9353: estado = 9354;
9354: estado = 9355;
9355: estado = 9356;
9356: estado = 9357;
9357: estado = 9358;
9358: estado = 9359;
9359: estado = 9360;
9360: estado = 9361;
9361: estado = 9362;
9362: estado = 9363;
9363: estado = 9364;
9364: estado = 9365;
9365: estado = 9366;
9366: estado = 9367;
9367: estado = 9368;
9368: estado = 9369;
9369: estado = 9370;
9370: estado = 9371;
9371: estado = 9372;
9372: estado = 9373;
9373: estado = 9374;
9374: estado = 9375;
9375: estado = 9376;
9376: estado = 9377;
9377: estado = 9378;
9378: estado = 9379;
9379: estado = 9380;
9380: estado = 9381;
9381: estado = 9382;
9382: estado = 9383;
9383: estado = 9384;
9384: estado = 9385;
9385: estado = 9386;
9386: estado = 9387;
9387: estado = 9388;
9388: estado = 9389;
9389: estado = 9390;
9390: estado = 9391;
9391: estado = 9392;
9392: estado = 9393;
9393: estado = 9394;
9394: estado = 9395;
9395: estado = 9396;
9396: estado = 9397;
9397: estado = 9398;
9398: estado = 9399;
9399: estado = 9400;
9400: estado = 9401;
9401: estado = 9402;
9402: estado = 9403;
9403: estado = 9404;
9404: estado = 9405;
9405: estado = 9406;
9406: estado = 9407;
9407: estado = 9408;
9408: estado = 9409;
9409: estado = 9410;
9410: estado = 9411;
9411: estado = 9412;
9412: estado = 9413;
9413: estado = 9414;
9414: estado = 9415;
9415: estado = 9416;
9416: estado = 9417;
9417: estado = 9418;
9418: estado = 9419;
9419: estado = 9420;
9420: estado = 9421;
9421: estado = 9422;
9422: estado = 9423;
9423: estado = 9424;
9424: estado = 9425;
9425: estado = 9426;
9426: estado = 9427;
9427: estado = 9428;
9428: estado = 9429;
9429: estado = 9430;
9430: estado = 9431;
9431: estado = 9432;
9432: estado = 9433;
9433: estado = 9434;
9434: estado = 9435;
9435: estado = 9436;
9436: estado = 9437;
9437: estado = 9438;
9438: estado = 9439;
9439: estado = 9440;
9440: estado = 9441;
9441: estado = 9442;
9442: estado = 9443;
9443: estado = 9444;
9444: estado = 9445;
9445: estado = 9446;
9446: estado = 9447;
9447: estado = 9448;
9448: estado = 9449;
9449: estado = 9450;
9450: estado = 9451;
9451: estado = 9452;
9452: estado = 9453;
9453: estado = 9454;
9454: estado = 9455;
9455: estado = 9456;
9456: estado = 9457;
9457: estado = 9458;
9458: estado = 9459;
9459: estado = 9460;
9460: estado = 9461;
9461: estado = 9462;
9462: estado = 9463;
9463: estado = 9464;
9464: estado = 9465;
9465: estado = 9466;
9466: estado = 9467;
9467: estado = 9468;
9468: estado = 9469;
9469: estado = 9470;
9470: estado = 9471;
9471: estado = 9472;
9472: estado = 9473;
9473: estado = 9474;
9474: estado = 9475;
9475: estado = 9476;
9476: estado = 9477;
9477: estado = 9478;
9478: estado = 9479;
9479: estado = 9480;
9480: estado = 9481;
9481: estado = 9482;
9482: estado = 9483;
9483: estado = 9484;
9484: estado = 9485;
9485: estado = 9486;
9486: estado = 9487;
9487: estado = 9488;
9488: estado = 9489;
9489: estado = 9490;
9490: estado = 9491;
9491: estado = 9492;
9492: estado = 9493;
9493: estado = 9494;
9494: estado = 9495;
9495: estado = 9496;
9496: estado = 9497;
9497: estado = 9498;
9498: estado = 9499;
9499: estado = 9500;
9500: estado = 9501;
9501: estado = 9502;
9502: estado = 9503;
9503: estado = 9504;
9504: estado = 9505;
9505: estado = 9506;
9506: estado = 9507;
9507: estado = 9508;
9508: estado = 9509;
9509: estado = 9510;
9510: estado = 9511;
9511: estado = 9512;
9512: estado = 9513;
9513: estado = 9514;
9514: estado = 9515;
9515: estado = 9516;
9516: estado = 9517;
9517: estado = 9518;
9518: estado = 9519;
9519: estado = 9520;
9520: estado = 9521;
9521: estado = 9522;
9522: estado = 9523;
9523: estado = 9524;
9524: estado = 9525;
9525: estado = 9526;
9526: estado = 9527;
9527: estado = 9528;
9528: estado = 9529;
9529: estado = 9530;
9530: estado = 9531;
9531: estado = 9532;
9532: estado = 9533;
9533: estado = 9534;
9534: estado = 9535;
9535: estado = 9536;
9536: estado = 9537;
9537: estado = 9538;
9538: estado = 9539;
9539: estado = 9540;
9540: estado = 9541;
9541: estado = 9542;
9542: estado = 9543;
9543: estado = 9544;
9544: estado = 9545;
9545: estado = 9546;
9546: estado = 9547;
9547: estado = 9548;
9548: estado = 9549;
9549: estado = 9550;
9550: estado = 9551;
9551: estado = 9552;
9552: estado = 9553;
9553: estado = 9554;
9554: estado = 9555;
9555: estado = 9556;
9556: estado = 9557;
9557: estado = 9558;
9558: estado = 9559;
9559: estado = 9560;
9560: estado = 9561;
9561: estado = 9562;
9562: estado = 9563;
9563: estado = 9564;
9564: estado = 9565;
9565: estado = 9566;
9566: estado = 9567;
9567: estado = 9568;
9568: estado = 9569;
9569: estado = 9570;
9570: estado = 9571;
9571: estado = 9572;
9572: estado = 9573;
9573: estado = 9574;
9574: estado = 9575;
9575: estado = 9576;
9576: estado = 9577;
9577: estado = 9578;
9578: estado = 9579;
9579: estado = 9580;
9580: estado = 9581;
9581: estado = 9582;
9582: estado = 9583;
9583: estado = 9584;
9584: estado = 9585;
9585: estado = 9586;
9586: estado = 9587;
9587: estado = 9588;
9588: estado = 9589;
9589: estado = 9590;
9590: estado = 9591;
9591: estado = 9592;
9592: estado = 9593;
9593: estado = 9594;
9594: estado = 9595;
9595: estado = 9596;
9596: estado = 9597;
9597: estado = 9598;
9598: estado = 9599;
9599: estado = 9600;
9600: estado = 9601;
9601: estado = 9602;
9602: estado = 9603;
9603: estado = 9604;
9604: estado = 9605;
9605: estado = 9606;
9606: estado = 9607;
9607: estado = 9608;
9608: estado = 9609;
9609: estado = 9610;
9610: estado = 9611;
9611: estado = 9612;
9612: estado = 9613;
9613: estado = 9614;
9614: estado = 9615;
9615: estado = 9616;
9616: estado = 9617;
9617: estado = 9618;
9618: estado = 9619;
9619: estado = 9620;
9620: estado = 9621;
9621: estado = 9622;
9622: estado = 9623;
9623: estado = 9624;
9624: estado = 9625;
9625: estado = 9626;
9626: estado = 9627;
9627: estado = 9628;
9628: estado = 9629;
9629: estado = 9630;
9630: estado = 9631;
9631: estado = 9632;
9632: estado = 9633;
9633: estado = 9634;
9634: estado = 9635;
9635: estado = 9636;
9636: estado = 9637;
9637: estado = 9638;
9638: estado = 9639;
9639: estado = 9640;
9640: estado = 9641;
9641: estado = 9642;
9642: estado = 9643;
9643: estado = 9644;
9644: estado = 9645;
9645: estado = 9646;
9646: estado = 9647;
9647: estado = 9648;
9648: estado = 9649;
9649: estado = 9650;
9650: estado = 9651;
9651: estado = 9652;
9652: estado = 9653;
9653: estado = 9654;
9654: estado = 9655;
9655: estado = 9656;
9656: estado = 9657;
9657: estado = 9658;
9658: estado = 9659;
9659: estado = 9660;
9660: estado = 9661;
9661: estado = 9662;
9662: estado = 9663;
9663: estado = 9664;
9664: estado = 9665;
9665: estado = 9666;
9666: estado = 9667;
9667: estado = 9668;
9668: estado = 9669;
9669: estado = 9670;
9670: estado = 9671;
9671: estado = 9672;
9672: estado = 9673;
9673: estado = 9674;
9674: estado = 9675;
9675: estado = 9676;
9676: estado = 9677;
9677: estado = 9678;
9678: estado = 9679;
9679: estado = 9680;
9680: estado = 9681;
9681: estado = 9682;
9682: estado = 9683;
9683: estado = 9684;
9684: estado = 9685;
9685: estado = 9686;
9686: estado = 9687;
9687: estado = 9688;
9688: estado = 9689;
9689: estado = 9690;
9690: estado = 9691;
9691: estado = 9692;
9692: estado = 9693;
9693: estado = 9694;
9694: estado = 9695;
9695: estado = 9696;
9696: estado = 9697;
9697: estado = 9698;
9698: estado = 9699;
9699: estado = 9700;
9700: estado = 9701;
9701: estado = 9702;
9702: estado = 9703;
9703: estado = 9704;
9704: estado = 9705;
9705: estado = 9706;
9706: estado = 9707;
9707: estado = 9708;
9708: estado = 9709;
9709: estado = 9710;
9710: estado = 9711;
9711: estado = 9712;
9712: estado = 9713;
9713: estado = 9714;
9714: estado = 9715;
9715: estado = 9716;
9716: estado = 9717;
9717: estado = 9718;
9718: estado = 9719;
9719: estado = 9720;
9720: estado = 9721;
9721: estado = 9722;
9722: estado = 9723;
9723: estado = 9724;
9724: estado = 9725;
9725: estado = 9726;
9726: estado = 9727;
9727: estado = 9728;
9728: estado = 9729;
9729: estado = 9730;
9730: estado = 9731;
9731: estado = 9732;
9732: estado = 9733;
9733: estado = 9734;
9734: estado = 9735;
9735: estado = 9736;
9736: estado = 9737;
9737: estado = 9738;
9738: estado = 9739;
9739: estado = 9740;
9740: estado = 9741;
9741: estado = 9742;
9742: estado = 9743;
9743: estado = 9744;
9744: estado = 9745;
9745: estado = 9746;
9746: estado = 9747;
9747: estado = 9748;
9748: estado = 9749;
9749: estado = 9750;
9750: estado = 9751;
9751: estado = 9752;
9752: estado = 9753;
9753: estado = 9754;
9754: estado = 9755;
9755: estado = 9756;
9756: estado = 9757;
9757: estado = 9758;
9758: estado = 9759;
9759: estado = 9760;
9760: estado = 9761;
9761: estado = 9762;
9762: estado = 9763;
9763: estado = 9764;
9764: estado = 9765;
9765: estado = 9766;
9766: estado = 9767;
9767: estado = 9768;
9768: estado = 9769;
9769: estado = 9770;
9770: estado = 9771;
9771: estado = 9772;
9772: estado = 9773;
9773: estado = 9774;
9774: estado = 9775;
9775: estado = 9776;
9776: estado = 9777;
9777: estado = 9778;
9778: estado = 9779;
9779: estado = 9780;
9780: estado = 9781;
9781: estado = 9782;
9782: estado = 9783;
9783: estado = 9784;
9784: estado = 9785;
9785: estado = 9786;
9786: estado = 9787;
9787: estado = 9788;
9788: estado = 9789;
9789: estado = 9790;
9790: estado = 9791;
9791: estado = 9792;
9792: estado = 9793;
9793: estado = 9794;
9794: estado = 9795;
9795: estado = 9796;
9796: estado = 9797;
9797: estado = 9798;
9798: estado = 9799;
9799: estado = 9800;
9800: estado = 9801;
9801: estado = 9802;
9802: estado = 9803;
9803: estado = 9804;
9804: estado = 9805;
9805: estado = 9806;
9806: estado = 9807;
9807: estado = 9808;
9808: estado = 9809;
9809: estado = 9810;
9810: estado = 9811;
9811: estado = 9812;
9812: estado = 9813;
9813: estado = 9814;
9814: estado = 9815;
9815: estado = 9816;
9816: estado = 9817;
9817: estado = 9818;
9818: estado = 9819;
9819: estado = 9820;
9820: estado = 9821;
9821: estado = 9822;
9822: estado = 9823;
9823: estado = 9824;
9824: estado = 9825;
9825: estado = 9826;
9826: estado = 9827;
9827: estado = 9828;
9828: estado = 9829;
9829: estado = 9830;
9830: estado = 9831;
9831: estado = 9832;
9832: estado = 9833;
9833: estado = 9834;
9834: estado = 9835;
9835: estado = 9836;
9836: estado = 9837;
9837: estado = 9838;
9838: estado = 9839;
9839: estado = 9840;
9840: estado = 9841;
9841: estado = 9842;
9842: estado = 9843;
9843: estado = 9844;
9844: estado = 9845;
9845: estado = 9846;
9846: estado = 9847;
9847: estado = 9848;
9848: estado = 9849;
9849: estado = 9850;
9850: estado = 9851;
9851: estado = 9852;
9852: estado = 9853;
9853: estado = 9854;
9854: estado = 9855;
9855: estado = 9856;
9856: estado = 9857;
9857: estado = 9858;
9858: estado = 9859;
9859: estado = 9860;
9860: estado = 9861;
9861: estado = 9862;
9862: estado = 9863;
9863: estado = 9864;
9864: estado = 9865;
9865: estado = 9866;
9866: estado = 9867;
9867: estado = 9868;
9868: estado = 9869;
9869: estado = 9870;
9870: estado = 9871;
9871: estado = 9872;
9872: estado = 9873;
9873: estado = 9874;
9874: estado = 9875;
9875: estado = 9876;
9876: estado = 9877;
9877: estado = 9878;
9878: estado = 9879;
9879: estado = 9880;
9880: estado = 9881;
9881: estado = 9882;
9882: estado = 9883;
9883: estado = 9884;
9884: estado = 9885;
9885: estado = 9886;
9886: estado = 9887;
9887: estado = 9888;
9888: estado = 9889;
9889: estado = 9890;
9890: estado = 9891;
9891: estado = 9892;
9892: estado = 9893;
9893: estado = 9894;
9894: estado = 9895;
9895: estado = 9896;
9896: estado = 9897;
9897: estado = 9898;
9898: estado = 9899;
9899: estado = 9900;
9900: estado = 9901;
9901: estado = 9902;
9902: estado = 9903;
9903: estado = 9904;
9904: estado = 9905;
9905: estado = 9906;
9906: estado = 9907;
9907: estado = 9908;
9908: estado = 9909;
9909: estado = 9910;
9910: estado = 9911;
9911: estado = 9912;
9912: estado = 9913;
9913: estado = 9914;
9914: estado = 9915;
9915: estado = 9916;
9916: estado = 9917;
9917: estado = 9918;
9918: estado = 9919;
9919: estado = 9920;
9920: estado = 9921;
9921: estado = 9922;
9922: estado = 9923;
9923: estado = 9924;
9924: estado = 9925;
9925: estado = 9926;
9926: estado = 9927;
9927: estado = 9928;
9928: estado = 9929;
9929: estado = 9930;
9930: estado = 9931;
9931: estado = 9932;
9932: estado = 9933;
9933: estado = 9934;
9934: estado = 9935;
9935: estado = 9936;
9936: estado = 9937;
9937: estado = 9938;
9938: estado = 9939;
9939: estado = 9940;
9940: estado = 9941;
9941: estado = 9942;
9942: estado = 9943;
9943: estado = 9944;
9944: estado = 9945;
9945: estado = 9946;
9946: estado = 9947;
9947: estado = 9948;
9948: estado = 9949;
9949: estado = 9950;
9950: estado = 9951;
9951: estado = 9952;
9952: estado = 9953;
9953: estado = 9954;
9954: estado = 9955;
9955: estado = 9956;
9956: estado = 9957;
9957: estado = 9958;
9958: estado = 9959;
9959: estado = 9960;
9960: estado = 9961;
9961: estado = 9962;
9962: estado = 9963;
9963: estado = 9964;
9964: estado = 9965;
9965: estado = 9966;
9966: estado = 9967;
9967: estado = 9968;
9968: estado = 9969;
9969: estado = 9970;
9970: estado = 9971;
9971: estado = 9972;
9972: estado = 9973;
9973: estado = 9974;
9974: estado = 9975;
9975: estado = 9976;
9976: estado = 9977;
9977: estado = 9978;
9978: estado = 9979;
9979: estado = 9980;
9980: estado = 9981;
9981: estado = 9982;
9982: estado = 9983;
9983: estado = 9984;
9984: estado = 9985;
9985: estado = 9986;
9986: estado = 9987;
9987: estado = 9988;
9988: estado = 9989;
9989: estado = 9990;
9990: estado = 9991;
9991: estado = 9992;
9992: estado = 9993;
9993: estado = 9994;
9994: estado = 9995;
9995: estado = 9996;
9996: estado = 9997;
9997: estado = 9998;
9998: estado = 9999;
				default:
					begin 
						estado = 0;
						clk_out = 0;
					end
			endcase*/
			estado = estado + 1;
			
			if (estado == 5000) begin 
				clk_out = 1;
			end	
			else if (estado == 10000) begin 
			   clk_out = 0;
				estado = 0;
			end
			
			
			
		end

endmodule 
module bios(write_clock, read_clock, reset, biosAddress, out);
	
	parameter DATA_WIDTH = 32;
	parameter BIOS_BITS = 9;
	localparam BIOS_SIZE = 2**BIOS_BITS; 
	
	input write_clock, read_clock, reset;
	input [DATA_WIDTH-1:0] biosAddress;
	output reg [DATA_WIDTH-1:0] out;
	
	
	reg [DATA_WIDTH-1:0] BIOS [BIOS_SIZE-1:0]; 			// BIOS_SIZE words of 32-bit memory
	
	localparam 	N0 = 8'h30, N1 = 8'h31, N2 = 8'h32, N3 = 8'h33, N4 = 8'h34, N5 = 8'h35, N6 = 8'h36,
					N7 = 8'h37, N8 = 8'h38, N9 = 8'h39,
					AA = 8'h41, BB = 8'h42, CC = 8'h43, DD = 8'h44, EE = 8'h45, FF = 8'h46, GG = 8'h47,
					HH = 8'h48, II = 8'h49, JJ = 8'h4A, KK = 8'h4B, LL = 8'h4C, MM = 8'h4D, NN = 8'h4E,
					OO = 8'h4F, PP = 8'h50, QQ = 8'h51, RR = 8'h52, SS = 8'h53, TT = 8'h54, UU = 8'h55,
					VV = 8'h56, WW = 8'h57, XX = 8'h58, YY = 8'h59, ZZ = 8'h5A,
					A  = 8'h61, B  = 8'h62, C  = 8'h63, D  = 8'h64, E  = 8'h65, F  = 8'h66, G  = 8'h67,
					H  = 8'h68, I  = 8'h69, J  = 8'h6A, K  = 8'h6B, L  = 8'h6C, M  = 8'h6D, N  = 8'h6E,
					O  = 8'h6F, P  = 8'h70, Q  = 8'h71, R  = 8'h72, S  = 8'h73, T  = 8'h74, U  = 8'h75,
					V  = 8'h76, W  = 8'h77, X  = 8'h78, Y  = 8'h79, Z  = 8'h7A,
					BLANK = 8'h20, PIPE = 8'h7C, EQUAL = 8'h3D, LTHAN = 8'h3C, GTHAN = 8'h3E,
					TIMES = 8'h2A, PLUS = 8'h2B, MINUS = 8'h2D, DIV = 8'h2F,
					QMARK = 8'h3F;
	
	localparam  P00 = 5'h00, P01 = 5'h01, P02 = 5'h02, P03 = 5'h03, P04 = 5'h04, P05 = 5'h05, 
					P06 = 5'h06, P07 = 5'h07, P08 = 5'h08, P09 = 5'h09, P0A = 5'h0A, P0B = 5'h0B, 
					P0C = 5'h0C, P0D = 5'h0D, P0E = 5'h0E, P0F = 5'h0F,
					P10 = 5'h10, P11 = 5'h11, P12 = 5'h12, P13 = 5'h13, P14 = 5'h14, P15 = 5'h15, 
					P16 = 5'h16, P17 = 5'h17, P18 = 5'h18, P19 = 5'h19, P1A = 5'h1A, P1B = 5'h1B, 
					P1C = 5'h1C, P1D = 5'h1D, P1E = 5'h1E, P1F = 5'h1F;
	
	
	always @ (posedge read_clock)
	begin
		
		out <= BIOS[biosAddress];
		
	end
		
		
	always @ (*)
	begin
		
		BIOS[0] <= 32'b000101_00000_00001_0000000000001010; // li 1 10
		BIOS[1] <= 32'b000101_00000_00010_0110000110101000; // li 2 25000  2 deslocado
		BIOS[2] <= 32'b000101_00000_00011_0110000110101000; // li 3 25000
		BIOS[3] <= 32'b000101_00000_00100_0000000000000000; // li 4 0 / so_begin
		BIOS[4] <= 32'b000101_00000_00101_0000101110110011; // li 5 2995 / so_end
		BIOS[5] <= 32'b000000_00010_00010_00000_00010_000000; // sll 2 2 2
		BIOS[6] <= 32'b000000_00011_00011_00000_00001_000000; // sll 3 3 1
		BIOS[7] <= 32'b00000000000000000000000000000000; //noop
		BIOS[8] <= 32'b00000000000000000000000000000000; //noop
		BIOS[9] <= 32'b00000000000000000000000000000000; //noop
		BIOS[10] <= 32'b00000000000000000000000000000000; //noop
		BIOS[11] <= 32'b00000000000000000000000000000000; //noop
		BIOS[12] <= 32'b00000000000000000000000000000000; //noop
		BIOS[13] <= 32'b00000000000000000000000000000000; //noop
		BIOS[14] <= 32'b00000000000000000000000000000000; //noop
		BIOS[15] <= 32'b00000000000000000000000000000000; //noop
		BIOS[16] <= {24'b100111_00001_00000_00000_000, BB}; // noop / _BIOS__STARTING_
		BIOS[17] <= {24'b100111_00010_00000_00000_000, II}; // noop
		BIOS[18] <= {24'b100111_00011_00000_00000_000, OO}; // noop
		BIOS[19] <= {24'b100111_00100_00000_00000_000, SS}; // noop
		BIOS[20] <= {24'b100111_00111_00000_00000_000, SS}; // noop
		BIOS[21] <= {24'b100111_01000_00000_00000_000, TT}; // noop
		BIOS[22] <= {24'b100111_01001_00000_00000_000, AA}; // noop
		BIOS[23] <= {24'b100111_01010_00000_00000_000, RR}; // noop
		BIOS[24] <= {24'b100111_01011_00000_00000_000, TT}; // noop
		BIOS[25] <= {24'b100111_01100_00000_00000_000, II}; // noop
		BIOS[26] <= {24'b100111_01101_00000_00000_000, NN}; // noop
		BIOS[27] <= {24'b100111_01110_00000_00000_000, GG}; // noop
		BIOS[28] <= 32'b000000_00010_01010_00000_00000_010000; // move 10 2
		BIOS[29] <= 32'b000000_01010_01010_00000_00001_000001; // srl 10 10 1
		BIOS[30] <= 32'b000101_00000_01011_0000000000000000; // li 11 0
		BIOS[31] <= 32'b000011_01011_01011_0000000000000001; // inc 11 / sleep1
		BIOS[32] <= 32'b001000_01011_01010_1111111111111111; // bne 11 10 sleep1
		BIOS[33] <= 32'b100110_00000000000000000000000000; // clear
		BIOS[34] <= {24'b100111_00001_00000_00000_000, SS}; // noop / _System_Loading_
		BIOS[35] <= {24'b100111_00010_00000_00000_000, Y}; // noop
		BIOS[36] <= {24'b100111_00011_00000_00000_000, S}; // noop
		BIOS[37] <= {24'b100111_00100_00000_00000_000, T}; // noop
		BIOS[38] <= {24'b100111_00101_00000_00000_000, E}; // noop
		BIOS[39] <= {24'b100111_00110_00000_00000_000, M}; // noop
		BIOS[40] <= {24'b100111_01000_00000_00000_000, LL}; // noop
		BIOS[41] <= {24'b100111_01001_00000_00000_000, O}; // noop
		BIOS[42] <= {24'b100111_01010_00000_00000_000, A}; // noop
		BIOS[43] <= {24'b100111_01011_00000_00000_000, D}; // noop
		BIOS[44] <= {24'b100111_01100_00000_00000_000, I}; // noop
		BIOS[45] <= {24'b100111_01101_00000_00000_000, N}; // noop
		BIOS[46] <= {24'b100111_01110_00000_00000_000, G}; // noop
		BIOS[47] <= 32'b000000_00011_01010_00000_00000_010000; // move 10 3
		BIOS[48] <= 32'b000000_01010_01010_00000_00001_000001; // srl 10 10 1
		BIOS[49] <= 32'b000101_00000_01011_0000000000000000; // li 11 0
		BIOS[50] <= 32'b000000_01011_01011_00000_00000_001001; // inc 11 / sleep2
		BIOS[51] <= 32'b001000_01011_01010_1111111111111111; // bne 11 10 sleep2
		BIOS[52] <= {24'b100111_10000_00000_00000_000, GTHAN}; // noop
		BIOS[53] <= {24'b100111_11111_00000_00000_000, LTHAN}; // noop
		BIOS[54] <= 32'b000000_00011_01010_00000_00000_010000; // move 10 3
		BIOS[55] <= 32'b000000_01010_01010_00000_00001_000001; // srl 10 10 1
		BIOS[56] <= 32'b000101_00000_01011_0000000000000000; // li 11 0
		BIOS[57] <= 32'b000000_01011_01011_00000_00000_001001; // inc 11 / sleep3
		BIOS[58] <= 32'b001000_01011_01010_1111111111111111; // bne 11 10 sleep3
		BIOS[59] <= {24'b100111_10010_00000_00000_000, GTHAN}; // noop
		BIOS[60] <= {24'b100111_11101_00000_00000_000, LTHAN}; // noop
		BIOS[61] <= 32'b000000_00011_01010_00000_00000_010000; // move 10 3
		BIOS[62] <= 32'b000000_01010_01010_00000_00001_000001; // srl 10 10 1
		BIOS[63] <= 32'b000101_00000_01011_0000000000000000; // li 11 0
		BIOS[64] <= 32'b000000_01011_01011_00000_00000_001001; // inc 11 / sleep4
		BIOS[65] <= 32'b001000_01011_01010_1111111111111111; // bne 11 10 sleep4
		BIOS[66] <= {24'b100111_10100_00000_00000_000, GTHAN}; // noop
		BIOS[67] <= {24'b100111_11011_00000_00000_000, LTHAN}; // noop 
		BIOS[68] <= 32'b000000_00011_01010_00000_00000_010000; // move 10 3
		BIOS[69] <= 32'b000000_01010_01010_00000_00001_000001; // srl 10 10 1
		BIOS[70] <= 32'b000101_00000_01011_0000000000000000; // li 11 0
		BIOS[71] <= 32'b000000_01011_01011_00000_00000_001001; // inc 11 / sleep5
		BIOS[72] <= 32'b001000_01011_01010_1111111111111111; // bne 11 10 sleep5
		BIOS[73] <= {24'b100111_10110_00000_00000_000, GTHAN}; // noop
		BIOS[74] <= {24'b100111_11001_00000_00000_000, LTHAN}; // noop 
		BIOS[75] <= 32'b000000_00011_01010_00000_00000_010000; // move 10 3
		BIOS[76] <= 32'b000000_01010_01010_00000_00001_000001; // srl 10 10 1
		BIOS[77] <= 32'b000101_00000_01011_0000000000000000; // li 11 0
		BIOS[78] <= 32'b000000_01011_01011_00000_00000_001001; // inc 11 / sleep6
		BIOS[79] <= 32'b001000_01011_01010_1111111111111111; // bne 11 10 sleep6
		BIOS[80] <= 32'b000000_00100_01010_00000_00000_010000; // move 10 4
		BIOS[81] <= 32'b000000_00101_01011_00000_00000_010000; // move 11 5
		BIOS[82] <= 32'b100011_00000_01010_01010_00000_000000; // hdtoinst / load_so
		BIOS[83] <= 32'b000000_01010_01010_00000_00000_001001; // inc 10 
		BIOS[84] <= 32'b001000_01010_01011_1111111111111110; // bne 10 11 load_so
		BIOS[85] <= 32'b100110_00000000000000000000000000; // noop / clear1
		BIOS[86] <= {24'b100111_00001_00000_00000_000, SS}; // noop / _System__loaded_
		BIOS[87] <= {24'b100111_00010_00000_00000_000, Y}; // noop
		BIOS[88] <= {24'b100111_00011_00000_00000_000, S}; // noop
		BIOS[89] <= {24'b100111_00100_00000_00000_000, T}; // noop
		BIOS[90] <= {24'b100111_00101_00000_00000_000, E}; // noop
		BIOS[91] <= {24'b100111_00110_00000_00000_000, M}; // noop
		BIOS[92] <= {24'b100111_01001_00000_00000_000, LL}; // noop
		BIOS[93] <= {24'b100111_01010_00000_00000_000, O}; // noop
		BIOS[94] <= {24'b100111_01011_00000_00000_000, A}; // noop
		BIOS[95] <= {24'b100111_01100_00000_00000_000, D}; // noop
		BIOS[96] <= {24'b100111_01101_00000_00000_000, E}; // noop
		BIOS[97] <= {24'b100111_01110_00000_00000_000, D}; // noop
		BIOS[98] <= {24'b100111_10000_00000_00000_000, E}; // noop / enter_zero_input
		BIOS[99] <= {24'b100111_10001_00000_00000_000, N}; // noop
		BIOS[100] <= {24'b100111_10010_00000_00000_000, T}; // noop
		BIOS[101] <= {24'b100111_10011_00000_00000_000, E}; // noop
		BIOS[102] <= {24'b100111_10100_00000_00000_000, R}; // noop
		BIOS[103] <= {24'b100111_10110_00000_00000_000, Z}; // noop
		BIOS[104] <= {24'b100111_10111_00000_00000_000, E}; // noop
		BIOS[105] <= {24'b100111_11000_00000_00000_000, R}; // noop
		BIOS[106] <= {24'b100111_11001_00000_00000_000, O}; // noop
		BIOS[107] <= {24'b100111_11011_00000_00000_000, I}; // noop
		BIOS[108] <= {24'b100111_11100_00000_00000_000, N}; // noop
		BIOS[109] <= {24'b100111_11101_00000_00000_000, P}; // noop
		BIOS[110] <= {24'b100111_11110_00000_00000_000, U}; // noop
		BIOS[111] <= {24'b100111_11111_00000_00000_000, T}; // noop
		BIOS[112] <= 32'b001001_00000_01100_0000000000000000; // in 12 / zero_input
		BIOS[113] <= 32'b000010_00000_01100_0000000000000000; // sw 12 $zero 0
		BIOS[114] <= 32'b000001_00000_01101_0000000000000000; // lw 13 $zero 0
		BIOS[115] <= 32'b001000_01101_00000_1111111111111101; // bne 13 $zero zero_input
		BIOS[116] <= 32'b00000000000000000000000000000000; //noop
		BIOS[117] <= 32'b00000000000000000000000000000000; //noop
		BIOS[118] <= 32'b00000000000000000000000000000000; //noop
		BIOS[119] <= 32'b00000000000000000000000000000000; //noop
		BIOS[120] <= 32'b00000000000000000000000000000000; //noop
		BIOS[121] <= 32'b00000000000000000000000000000000; //noop
		BIOS[122] <= 32'b00000000000000000000000000000000; //noop
		BIOS[123] <= 32'b00000000000000000000000000000000; //noop
		BIOS[124] <= 32'b100110_00000000000000000000000000; // noop / clear2
		BIOS[125] <= {24'b100111_00011_00000_00000_000, WW}; // noop / ___Welcome_to___
		BIOS[126] <= {24'b100111_00100_00000_00000_000, E}; // noop
		BIOS[127] <= {24'b100111_00101_00000_00000_000, L}; // noop
		BIOS[128] <= {24'b100111_00110_00000_00000_000, C}; // noop
		BIOS[129] <= {24'b100111_00111_00000_00000_000, O}; // noop
		BIOS[130] <= {24'b100111_01000_00000_00000_000, M}; // noop
		BIOS[131] <= {24'b100111_01001_00000_00000_000, E}; // noop
		BIOS[132] <= {24'b100111_01011_00000_00000_000, T}; // noop
		BIOS[133] <= {24'b100111_01100_00000_00000_000, O}; // noop
		BIOS[134] <= {24'b100111_10001_00000_00000_000, I}; // noop / _iloop32_system_
		BIOS[135] <= {24'b100111_10010_00000_00000_000, L}; // noop
		BIOS[136] <= {24'b100111_10011_00000_00000_000, O}; // noop
		BIOS[137] <= {24'b100111_10100_00000_00000_000, O}; // noop
		BIOS[138] <= {24'b100111_10101_00000_00000_000, P}; // noop
		BIOS[139] <= {24'b100111_10110_00000_00000_000, N3}; // noop
		BIOS[140] <= {24'b100111_10111_00000_00000_000, N2}; // noop
		BIOS[141] <= {24'b100111_11001_00000_00000_000, S}; // noop
		BIOS[142] <= {24'b100111_11010_00000_00000_000, Y}; // noop
		BIOS[143] <= {24'b100111_11011_00000_00000_000, S}; // noop
		BIOS[144] <= {24'b100111_11100_00000_00000_000, T}; // noop
		BIOS[145] <= {24'b100111_11101_00000_00000_000, E}; // noop
		BIOS[146] <= {24'b100111_11110_00000_00000_000, M}; // noop
		BIOS[147] <= 32'b000000_00010_01010_00000_00000_010000; // move 10 2
		BIOS[148] <= 32'b000000_01010_01010_00000_00001_000001; // srl 10 10 1
		BIOS[149] <= 32'b000101_00000_01011_0000000000000000; // li 11 0
		BIOS[150] <= 32'b000000_01011_01011_00000_00000_001001; // inc 11 / sleep7
		BIOS[151] <= 32'b001000_01011_01010_1111111111111111; // bne 11 10 sleep7
		BIOS[152] <= 32'b000101_00000_00001_0000000000000000; // li 1 0
		BIOS[153] <= 32'b000101_00000_00010_0000000000000000; // li 2 0
		BIOS[154] <= 32'b000101_00000_00011_0000000000000000; // li 3 0
		BIOS[155] <= 32'b000101_00000_00100_0000000000000000; // li 4 0
		BIOS[156] <= 32'b000101_00000_00101_0000000000000000; // li 5 0
		BIOS[157] <= 32'b000101_00000_00110_0000000000000000; // li 6 0
		BIOS[158] <= 32'b000101_00000_00111_0000000000000000; // li 7 0
		BIOS[159] <= 32'b000101_00000_01000_0000000000000000; // li 8 0
		BIOS[160] <= 32'b000101_00000_01001_0000000000000000; // li 9 0
		BIOS[161] <= 32'b000101_00000_01010_0000000000000000; // li 10 0
		BIOS[162] <= 32'b000101_00000_01011_0000000000000000; // li 11 0
		BIOS[163] <= 32'b000101_00000_01100_0000000000000000; // li 12 0
		BIOS[164] <= 32'b000101_00000_01101_0000000000000000; // li 13 0
		BIOS[165] <= 32'b000101_00000_01110_0000000000000000; // li 14 0
		BIOS[166] <= 32'b000101_00000_01111_0000000000000000; // li 15 0
		BIOS[167] <= 32'b000101_00000_10000_0000000000000000; // li 16 0
		BIOS[168] <= 32'b000101_00000_10001_0000000000000000; // li 17 0
		BIOS[169] <= 32'b000101_00000_10010_0000000000000000; // li 18 0
		BIOS[170] <= 32'b000101_00000_10011_0000000000000000; // li 19 0
		BIOS[171] <= 32'b000101_00000_10100_0000000000000000; // li 20 0
		BIOS[172] <= 32'b000101_00000_10101_0000000000000000; // li 21 0
		BIOS[173] <= 32'b000101_00000_10110_0000000000000000; // li 22 0
		BIOS[174] <= 32'b000101_00000_10111_0000000000000000; // li 23 0
		BIOS[175] <= 32'b000101_00000_11000_0000000000000000; // li 24 0
		BIOS[176] <= 32'b000101_00000_11001_0000000000000000; // li 25 0
		BIOS[177] <= 32'b000101_00000_11010_0000000000000000; // li 26 0
		BIOS[178] <= 32'b000101_00000_11011_0000000000000000; // li 27 0
		BIOS[179] <= 32'b000101_00000_11100_0000000000000000; // li 28 0
		BIOS[180] <= 32'b000101_00000_11101_0000000000000000; // li 29 0
		BIOS[181] <= 32'b000101_00000_11110_0000000000000000; // li 30 0
		BIOS[182] <= 32'b000101_00000_11111_0000000000000000; // li 31 0
		BIOS[183] <= 32'b100010_00000000000000000000000000; // upmem
	end

	

	
endmodule
